`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Eiho2wIY+0yBr0uzSznxrrYb/fsVAyjGuXlZ85zykkIbNwM9Vrakib/UdqcFKXyi
lMjtqRvQnvRm3yOxJMsPtTNNnX1H4OJMv1xIfvNeU7Bwc9wD0Z749NO5VbYEC7dI
fxjBnnIjq/0LT3ivX5sG9i752LnmeYafIAidvxGlZR9bjXjEImbbpaV+HQ2O8aWs
7ara5SYiqm12xyaSD3dfv+s/rQyt62TzO9oVRDP0aOJhoDqVYcK51zhqgF1bV4QC
agN1oIkZl7fxspBeULyoCPYmf94dgQcmkY3Im3JuhRFWlIAc/2HQJ1iGV4O6oLWU
R64mC25XJGEB1YQZGSs8NQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
UcK6hRXrNEJ6tyIhZu87lE++xksHDFFigcymzVV+K/LiRiyq9vwPwLIZLjz83TUt
N6MiAAmk+LwZSxwVJiooyDky3kXHkW6zaK+wBjfxjKYn45VsKJF+PlfWIEiBrRuF
7ro9v9lFLW0Pld4U3gg51f62Vzso0Lfi3owNwoomzNs=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 78560 )
`protect data_block
GnC/2mmLzYnWTLq+jgYtJhGh64ljvctbrEvJbGZ0zQmejVY26zMtlut42/u//xoH
KdHYbq+2sCN5IEyhnlmldwetXNKfPmT+D6T8/oUFPh/hlMm0TBzoMux5Fbm1WmyA
32rtQ2kTqVFX1m6DbwX77PZnhWO6nP5QVR8tcH7bad5Z0QKAhuJaB2T81QRWYdJO
D4+oqftffkNKxEPUWqTWH+BEPT6o8WNzFxcyNImG69HLktWGRxUZkdVIZTXBsjXJ
13wtDcru5qIoj8Ap6U6DP1MVaAsMrCL7ItZo7oMZMKDA91a0r1TY+vkZarDVMkLi
YN3FccRT7igsRzT1B2s6CldSBZofQ5cytfCBxoUiGwM2YN6NzNCZpXl6eBoNiACY
BiKb9ost3acd+NtKzA8GP7K1WgCX6vsbFMRKnFqyeRmuSA+hxTSSrnh+x59WyOl/
PSmKxhsJ6zPr7uxIvHNxrq+39bCqa3gyaH2NdQzrepEBiPRPp8q8gjRvkmNSpag3
T1kRjuFFz6pR0VHZcM9EdwmOlOyEDmrn27/jchnY2X+s2FEJMzXUsuEtIvJfTDDA
iS8Qo+4/EKQ5UJdckhe1edMLngedRUAgcnwU2HNg9tVzRjvAM5l7axJRrSl66QyO
3L1/Gkh3AvjIXMuvoSkooaalWDCVEteLrIvfGI1JVAbbifIRIcYA0LB7KJRFYDVA
bHFhp7V1q2QzIT2WGSx1xTXkixrXZKQ/fYDVE4OH0XMeSZbRHzr+Mc1/Ni+tlPSj
Yrt0lcWTfF+W86Uad+jwmGdFV6/wHzepl3ASEXwqwS8K/mFOaQo17czdulEP8fu8
z3s4qvHNDM82F0elHl+WHYWfK23Z7q0NodOqKeRR/NM83p+jJgVrb2bFtCnOdOkL
7myLQq38E1XmfRWf+vvIqFGqkman2GajR5qSeVOFGLnjNDEHFfmY64tPv2q1KcN1
yfNUPtQ16y9+4epLnbcqX9dOUSyUarTRLBVcCwmXpALBau0asExuNvyD2MlE9Bog
y+Q3+babPETw+zLyIEp7jBBHjkAVrjtYXiTbF76puaZ+nTuWvXVcqQ7wvfNhCE3V
veAet9fATswQc+RQWufcLAywm3Dbvd3NFBX40fgoF8gm+t67Zg4a7T7OoX8RVR8T
7leZY2G0nMPvO/B2cehddSCPlAaBhR1qUdj1y/Mrm5GetLZrH6J1Ps9n4t9Pyo/R
UAx47v+q+e+wncRdJcOxeHODMYbNy2MBpCHA/fGeHPMJUNpR+pgn5YH4uX/dPWMo
73ideqowO+xtdkJhJqaYGePG+2R2V542W3q2HqrZAtfavJRIp0yqJqraJRrxPgsp
KldMXBvdEGUpF9neRTG5eSGC2kKlenhbIX5YoenoQ2ExY9OMMv5QnugWP7WQlzjd
BWlQdTJyF36rLcaDeXhXrLCbuV/6fQA65+RUixopbVZarE1dnbRUyUcr5/k6QEsD
Ie2NTtuPWGAKSG6DWTeN3qizYkGGXZ48rA2ojrJUi929vcowS8iBkYqs19WAwj+T
QJkZFVtbvVfXCd71b2qlFX12CvWtoJT3PEAp7kScYCfXTvIJUKgodvVlK4oWeVp5
PG1e5/v27ZtUOirW6Jbje1ipUZs1QDB5UVgDdHE7IxRUEC5Tx4k138w9zO+UBop2
WecZO8jFEKVLEhLlSbeTAkz1S0njYJy2TbzPmSi/uiR4Ss31aKhtrDbaeJfx5Sg9
uPPlKlJD7jaCq+ec865nVefGWOPgsHkkeUTasF0lCOJfQD7JnDLYAFZN0DuVQYAQ
/SOmYnF9hECwAR6FGNOZCbrRPrdoJwH66n79aRp8xuMoPC1xkbFg66YJyeOvww/f
aF1Ww5qX828Id0KEDs9mqe36vI9QPKqE4EfbAyaTWiA/LusxFm0S+a+SaG/rSl5o
WDi5R+OUjWvBZxdYBYQYpAA4LiX1zwhh3MrzHvtAbZWbz+W43HYSOv5FlSqfY2oj
CvVStlYcwyr7JCsRBC9uBJuQWnKcnW8gG0jfgp3Dx1E+Liyr9LP3dF+wruhS6zAl
hzdidppK/xNw5+atFNGrayzd5PbsU9qvqQ9ZDeuDP1uaR3sshEiMxiJbbVNfi69J
TQfQenHCLiHtHmpPmtlrjplLbET/TTUoKmaB0n4BOGQra/grIIVRohFTQW7mbgxK
HYYaYUkkvsdTfk1aGoeB1o91HU3AopPtTwjKdlMaYtHb9WyQQvvMlFllJHJehTeA
n+Qj6hsjmwc7KHtEI4lvpbC/dXSLvSbg2K9X6TZv+pEo+0EQOvswtAlKSKgFflK1
nzeGZVWBVJoW+O41PHsOnyFYb06UTN70nAK32D1kSO6KzhhRL0S+S03N6EeSu7pT
K0U1BjiywgZDKSZlPfc99R1MMDW3TKmcgY7f8+G5eEkHFVhQwoQxKld+F6XTw1Dk
8kcre2p3r/Tlq4t/bUXvA4oBhOTn1zwAMiMhEpoyQdSypMHVjP5TkLrkeVR1CIfZ
S1XxkbfaWUdGpKxs0prJIvrcHXhkHvS0LoD9QNazr2NEbpsRneNaQhViedrDsT1f
2kau3LLkQc6hBzk3tlokRY9ZBDrU1ZsGQVJ8TAjoVCzgFw14TYQEMAy5XVQYlTff
/S8rE8Ar9M1XRGnSqKXvzucIhWoAwa6OM+I0d3J8EE9/AougQxh1vI6mx+/Mt5O4
QRTsRaolB6l8kbudzkej6RH5cdg02qJ4A9bxiUROy6t2O8W5HcgyL2JE4GSDe4Lb
Oj0GNkWkjxzUydL9Qc+/Dubt7tJ/gibLxZn129uS0HlV12sM5Monm2OXZ0XgxYl9
DYSbNMrj5pbf8gVIOYT6cugH0RCpbzXfDOMo4hJsOgIuxkbc+EXv8cfwOgyqbXWe
o8ZwS1OfD9VIj3UpJk3ebXNJ7WXys8n0UyEmoCRPEr1u0G6TOTxqqgG/UT+oU91D
uhklU5dWHbHfDxqCIsiGMuOBfUT8wLgWUXDx6MFGv1UcaSIchuUYWK1uCu4WQOKI
KntriMZUOchbTV4W1ddejmgVkoeZ+7J87PRl2N9cotu7uw9zv7Wtj5fA1zRJQL4f
TuErOvUYQ172tEdpWk7o7rGkRvKFKHWY2adwJqOTtGw/65vHRyXIRUPB39WN+jY+
BgJopSjYLlm2ybo323keFfHJahaRSMN59pZrhLw8fAS4ct3ROKclEMVcDEUZkP9J
2x7Waa8Pwy8pcUumblwI6GYGhhhElw5cV/5a7XDqHJD5l2oOiEW5jJjlPP90f8WT
FaATxTUAFOS9lc7veKG2RuWmS4pGt+SmfHdoVsUblxQwPKSxzWERSNdxVXpeeLxt
YEPtws9OpSoZlhMrSj/JQv4//kQfRgWoTiguZF0VHMSFSpw9XYt0go1u3YSYMhKT
F8zeGYtIrHwBsIQKbobVPFFwI8PnvwaMAhTshSLEwMrmrfKxqYRoH1/usY0qKDNI
uEzORfkuRC9qxwfk7R5WG0AnX4Dhml+Vx/UtWGKx3DQ06ZGm852Mukvb0HK8flPX
S+TBF/JCyibYZVTK5HJlPrWUBZDoWKggYg6NH9YqUw0LrZkaFycvJR7NuQkY/Msg
tF7//xQQiSEQ0wbODFN9dDNnF40tKD8kfTvOWXDVeCSEs7gv4JuThKZjOlfE6Laq
UIQhD+sACOdCzSx6HqU7WO96SG9QkQHdnpm1TokNzHFPzX5qdD59I80CO45+5dJF
i1ejfLQiwb8UTenPn95AK0pjAR9wZFGMlHD9yPRrWwIaY6F7P7US+kLwcOyq0J54
6+25DGJSap29nIxMJv+1Z/NzTpM6sjAmSL+WSkyjQIxT9yhpblS2qyl4uWa7oanR
x1WGRsDTao/yGVI3ZfvyFCfmvnL1uZTJ+rkeklFAFQ0b+J+u20Hez9xfti/v64o2
Wvnyy3aXf1+XIPYjK84B6evZv7l8kUf42UBMRI4v0YLRx37eSl41R40IU1yE92FS
yALtQv4qhoAJCtYVMw5RX0knWJVVJ7/WmYcmypRqGGvaQCmbxZDSaZklDzOm8cnN
dLNy3NQr7BM2V0p+yRYRyyWXRQHO01Nqklol5cCq3Ve3f4o/ul9vwnOQIYBBo34r
/yLMfM0bIlN0gFF8xAEtLPHbzf/nTALTn7v4xs7PjyBB+JBnJGoiFVZn/m2wB0+R
DIouJw8jUlEO5gTc66LdWazrhC67NeUN6EHTbtimMs0+09WetCbRzDSwL/XeIgfz
80pjt1en1wAB5kfdbeYT0xmX2J/FtLSxU60CHROc8sC8DrITNkfDO8F2RxFt91O+
nDBo//hUYirrC1Yky4LPb+GA/zLmCmuovcSq9e5rMmN7pT9DEd1qKPFNuvQeeJks
koOGLUtbTrPlCsLREtnnk5jVSk/JX9cpbpw4w9uJze0IXJ5ea7gzu+ciPuE24l85
tpdJUldcjFreksWOMpfoaB0nkux+qmlbe/laEX9Hg1S6irlQJtgHm02NvbAv5/jX
U6x57oG3UIqzhSLT6xPuGW9kai4kVvZ1T/0u/eOEACewxwWFa0tIHss0SEpe672h
5ROMKWCforwXiVM/uF732lfbpEx+aHEy2sQU37xf1WQFOye+L9iraksrYGmKNWkW
3nnYx7tAvAmZGiAYpSZjofyKmySKm12D/QNZgWSAVmWSUDFwNuhDjMGp1uts7kb5
AROxEFxnqZqv9fpiHGttoMVJn6kfX2rt1dT3F+44WqZQE9rJXrNkBZFR/EsSXWq/
ITebFQ10eS99iGohiPxKFqGemQifam5hfvF62K+BPHpO4Cd1s0Wz348QvgVnm0SS
hXlwaEICcJFH6uEdTyzakFf9nLk9zQHvw7FdKJ1B3I19NHMWfNTLHcYzv1Tnp68z
GllII9WEvvFq/KdQwnbMRqAUASTrTlvB+7u9Ljg/6YCbLYhUcN4v0jVdk2fi+NMB
OuoAX7/wg+mNa/wNCRQhvfuR+qugErKwkwQ8Cga60qY+fGMJTVFT34fROP0HLgRE
TGzYSDpCbnxeeGN1g1WJUlBGLvjaYxTXA1gx3bEPWBWD/EdBWD8AdQYAonyceWAn
ykzMwVpbG0JIHoI7rR44Hfjw/yHTKEuX3LHVxUB3GOP9yQDEo+rEk4GTPha3CbNx
vc27qLOkZpsS3ZNFqJ5pBK4OsHi4ufBMUW/dllRS/9Kcj+qxGqh8QC9OK8PV7HWs
SjPn8d8acorPxV28Lc3KdCK29y1ePrV+pQk7MkZl41DPHM0l/cGAofGYJNkKiY0z
GU/YACklkB2eHu7IaXgcDFdAl9qIjmrX22Yn0toaTue934baWZBmk1NGtqMN9JoS
Yua/sQcAihfDhYZqVDwUHOmQvVadPreLt/vY8LGh/g4nFIEzkW7ekgMh1tVP/NGQ
Vjb+rnOkFhjgyDn0YLQStMrSet8X0HWlojB1WnlGfJrcFEI2zoc7DRQsq4hO/7zG
dFgMVYnw1FoqaZmLS9hshyNtyVK0r+w8Dz3AC2tOWJNNmyXmWN2e71DWQykpkcWk
RREwnK0vmXQ9dzh0LYJzbwQqqPIP3q5IRgzjoVO6Exb3vF4AQRDFdZsSaxwQDuzR
Cz2QkkUZ6pthHxETbFdUZH2P8XYviUvmm+xcqJJElGYrmQdv3sSE/+qHdqZCFkB7
MxTVnQ28yeUtRp8EKCcId1cBqEnLxHAy/lWQ8555ACZwBR5cts3TOooeHdAcd+sd
1n62PDE5JPfnc30WSJcZr2GcNvP2lyWgDH5QNKfoFDXWytVIybuUAetLhYD00JGG
9BMkpJu6uWvQOgmpqivritJqQOIf5vX9qorZEeOfYpj5ndxzx0soRf5St/Ilwe1+
yUrSpuyWZlUXQQ2OcdtglmMkvwDQ6mm264P92XVoA+RcRcEsK2QA7zMNBR1Xvm3/
vLGtvvGESbJHp2VEhJvomETYAGWX77alGkDUYbsxi4X98f8iLjOG7u+yEawWYu37
yq1KX3lYRPxOWZ7j+VNQeBx7hUclRjcw/3KtqCPfbnK4qBthZd8YPr8U2VdcoLBr
0l4E21YhYlckqjCwAbiOWvICw1fPhLi4enevIJ3Azk4KvZYiuIhETc5y1Ydf4GkK
3CoaueWv1C68pcymzM90cJgvUlCpeWupmcadheHLWfP2PqRAU68VcxrNDJU6Sq26
/lrFXzIhkxDNaJ8HpXDB5QJLfGMjFUYjEVVaooVu0f7ijuCnFXvNLXz4xpsm6UIg
hfqeKRnyxnaAiCBw59xjcQoFZ/ImRDkE8mkmXAOgjUdopyGkeA1swwS8COSS44xt
6PAA4j7+jHVleGfaNr4grQJfD6W76sL5mqJ8z065BHaeALQ4I2derCupaw23yN+5
8ZD7N12BTG8oxHLphnzgUoolwdf2GvF0Vhc24/dL8UpuEpjmD9I/ASGOy1L/MdSf
fMsyMjH9GgINf2BOIeHUv+28GCimCwF4bboRlJi5m5csRYxMNh/2UZKg/9Y5lkRJ
plcTYZhQjWMj/atMhlUE/CjeM23mny3qZxKGSCsIAlDATJHZ5+oKXXD/QYNO2C1i
wuHPhumntocvF/YyZdtSTWSQZqYT0rhOswmCnjQKaJnYRJ5m/M4SN5+SBv+lMlQo
p1ZQflDzSd58EzEVnd1jfFDPulGBXRvLkZv5DnTQc54HRtG55volWxALdYZ9xZgg
8JAWAn6l4UfyzhqZNB/odrwJN+IDUno0p6uukE17hSnxJHzvtM0p11dqXeE0DFvh
t7dp9KGo+GVUYt5Hs586G9cioQ/jTq1WrMH5GE0V84XLbEvCf47Kz5BG8bpwGdS5
pPYMiR7vktk5wHAqOJaa/Nd059XQIwwef7aTomahrcGuozF8fqR2Zv8mUEtuFZys
NEx08OZSYzA2YSpp7mH5xDRfhBsEpz4v0wzlZ4W3W0/tzlSEvf1ldY4Gxc1vQOul
LHqUJT7SfMhfNqtVfBdocigmIUA/Gbv3IkIbRJl70UMxR3gj/Xk98bkywul0CPjl
dVrPtWLO1whnEFdmCWxmQ3jCplYlrsri/vb+cnDjAte2e1LYd2nq6S4md4VN29/n
U9ilVq28Ra088SqDSCzInqYabKQpf5fMB2sTEleIdE5QxsD6Wrqdk0oTWJRGPSju
MUbMs48BNfA/yWAsJIjOruDeF42vUhu5PrBhXzBWOvIlczn5s8cYBIhueqsIYJwN
S57taFLSf+oJlkDhB0M/PEfstiLG4K4QT/a60amUGUvnLmtgxaM0wB5+RZ2Qjlma
vspONP+Nzds03ox6PVRqf4Nyz58D+zx7n/jNxuYwAYqalSxd3GZCTLx7YT+o8xZw
Wq6cdDu4Q46//2EuDwiMMedwkV8AFw/HPxuXEPkzyGO85ie9sK4qw8OedBCk0/Ne
oDl01UjLSQ60tcZwoysUo/ip/TTkd1BIF2txa4mVBbAwETVEQSwsp9/KFMAZmOkm
woY4Pd8gpFspY+Vf15qodjLqCsQCluQWDLAqGveE/3ScdOrSjhG8NoW8jv3uxNax
SWvPir38/sWDL/1DMOVAunbPj9aEJnkzyF3DOUfzPyxR0gnFc7yBCeKcfGfI1+Oc
RMHrd1BTpu/qRkhHSi0qoR9RvVOFqT9GwKBvjMQ3HzF5GJWjtcTPxi/zLuR0BbQn
aNxvIv18VvuDztZTkzyguggzMKMYPH6MCoEm6MxUEGLvFPUIH5blu0CBItupwIDs
GOy0CEjTVk26HyAtYeL1kfgoz9Hp4EtaQ0OH3OyinPxxMWaF3kj+kzUmzK4+XgR1
ts0Phc++dicq/5HhAfFAWxDF8eUzs6Qs1daYv5PgShO7uF03M2CTp2OryeZ0+gAk
MQ2SFHUwLbEE6x0NwvjWNY5fbnO4k+5IcPfkGNth/V+d8hHv8RpDbgZlIMevWkIH
QCWnCjSs4URipnjudeusqo5+m/XEs/Wv5jCb3r5O4TvgNWu0fraJiFNqFkyA7Tmx
FSj3AK3vb80j0zitv/tggkFJ4wGuPuSjTUQqgCUBGKx74ztCYAFBAZbillUxauep
KPLUCy6H4AJ+IlqCEFj6fy1C/N7S8L0Bqips3PssfVY3non2dcb/7aj55kJpLfKz
8H042vJMBnQI5BvCM5BvC0kTK3XwecaQ9GwR35+aCiv55h/n60izq7hiMr9L7GCB
Tktk+iGqR/ToYT6uYdhOfySzgDmVSkYlgrgfl4B+msAVMZyqW4YP4l9Ur0hV07bf
JwO4rvTZJvHHRZMlkX8QehE3CVLinrv0PHu6LYA5elRnCtOike1K6X73SwcnemZ6
dyFepHwDPwEYX+lG779ERLQUpeiFwxAJtEPSr+VmzeL0PuFid/mWVhEE/UY17fOp
zuVqv8khssoYtBKYCYZTcPNKuBXqzu/3NXruFxBwbFdF8RmNXglvDqowebf7bkgo
ZkHTu/cNaH0nevqTsOerzdI/w/OxMQG4++S3OWdWAG5keytSmRpL1cpyh9MGgFCc
iftQssnMwdqSYqHq0BM/8JZqFbtCkIO1DtZVcRU16rMtmxgbOn8G0yfqZiuJCwXM
LHPcF3wyjA7lGZEKMjt9j06r/9DT8vcZPXasmvFLN1/86QDsQLPNbxzT6BKrpZnS
mrG5Tn4pqn6uRpfUx2JYNDVQ4GpW/RRghV8+RwFcScaj3h2vanmRp8i2uC1c+Y4P
1NdRL9q2z/Ty4pKR/fJkqiT7H04BcLR5cFayxWCAvMLDmtjm+QHD9D0oQxcOja1r
IzlKbu1H55O5H/TiDRYjiqAQXdP6rc/poCy3+Zr21CRZTUrjxuY8bupnCsEA3BMl
OXk4kPStz2gdoj63n8lH/UlO2s5YcdxUSLsAF+LsJAXEwccwj3Rfn/2YB7w5gVgj
EevVlMV5cSfOogQDWpF6csclUBneCrxrj47uUZQVQXavza3ha5uo1AUY/gB3c4OY
46nBdraDQzQwfyjTFnGpXQUBJ/3TCNMRXlxpzrIc/AzC/RL7yghXXuF5DGsVVOUr
HJ5sdobPKHtQrgMzcgN//Vrpp6OeVTuXMISeBXE/DIn757y6SL84FJQCVxmps91l
9bJ57kiy90zz8S0zdT4dUnmpiNC21n16tBPSwsDkQ2g/fQhWQlg+6TUi3464LoIa
p0bKHb1o+b5xX63D5AwER2SE+Sp0fy6y5TDjU+yQCHsHOXP+BmuGIPU7Pc6Nx18x
qNy8IFFLht0GRwTL3Aj0fu/9o2YWKkLGOanEG9K5oRGVEviCfHdCE38BDHYLh2ZR
NTZHWthiHAx+JlgX1YmgAH93UxqnYWI+lcLZjKC9aYNCippHYuZRASutVMbBRasU
3Z0PVUTli6LlIuoAPo2kYJO9TUwMBPv906AbcsFqk3AgHJ8lKlr2G3CyNMz3XtlD
E3pdwc7U0X5S9O7IjRPiD7SWtgF3Z5732BJqKPwd8Mge/8IPc/EAq1woUazbpZFG
k+7mg0lKa9P7MesoCR7f6spSbMGfy1kn6fhztCve4tcmBR6TvlpWfh5SJ87uYbOj
raoZWlvIB+lxsIb52tljCqvrGbcLjBym++jbi0mT83kmzoffdjcXRhrJprQgZz4f
oMcHLG1zee3WAoDZx9oN21IyI2LVt4crjlBOHLV//D7gEmCopuG2U6wGaNYmw3ho
CK1/WPwIliYDkstAiQf4NqppI8rat4b/mmR+5Rkm4kQpFOm22ODo3KkCWsVPORnD
u1fo3k5i1XeCRyoYZ3ExrTRob+GgfX/tc6Qv+0KgfAX2TO/IvE0BgDJio5Ca4xFl
P0Y238gYdQ42IkRBhlkrT+ohD+0nreKj2U+Jgp1YL+ep+9Ch5T9oipImOuklyaOw
O1kEYT5ZqQPDTOnY2jQVZzrUGoPfydxUbg2wqEj37yD1rAEvPcIaPa6CUJ63zqLy
5kr8xVQZiXs8uNA2wlp91BvWnLRsfMXsG0vR9zSg8h6GknEt5RBmdglBtXeb2+9g
FGkikqdMrjz/CTgdOgJ3CdT+nP3dVli+RumCN6SrvDALlF8ynq0FjdK7Ej69bwVa
BwJILEv81HK+uNTHX9BbismouRbgoEXoBYagbcIuygD4nVFKZ5rx+jRhE9GJTVwO
fuO/zu6kkJ1BcaHuDxPJaYNpedeeHl+MB88Od/SFlNr1i5f7No1KtJrwHo6M5/8p
d8WOdNhrdg0zWHuaQDe0u6Z4/nYV/73LJjJiek4yIjPmwuXxoEorNBgJfu2IfR+U
04RlrjQYpXOoIRLLzsT2Nv54vfgPI34we6vLJXwi3pbGa+q4UxzZreksg2N2EjC3
Iefykn6J66BYe4z2R7nTmEQuYLaAFQdVAeHlSfZfBY0ggJCol9oEcPybJpkvebCd
qaVdyN2WbdzhPLMXhUSNGuaXLh1rOl0F0uL+eshWgMNruH2sP8M2eKE2XMKeM1h2
TlMFwBLsqTziDPkkBygT7oUWm0FDCsiHQqz4rSLykbQy2Tbxfkzivud1mAJs/M5F
qP/d5nJXZAdw5VUJITWQFkOClSIyG7+nnk1NATaJ7McPBVOSwh8LXBYSnO8hxudy
Wjs1y26Vn/G6Cdq2u0rM1fK1JTFj58jGbxuKxbfqoXuCZWUaie8HnNcRpea2R/yw
t02sVezMZWLX2OjC/9a/bodOCtLFHICYBSOIHAEsdFuE2hkobIXs547SIxpeh6yY
TVdx6kNvwKb8yKankzAxO2Nfk3DL4/9R2z4d+F0hTDywPBdn03PqrRxsnnHvG4jh
J/C2eHc3fNnZCib1+2TXk2spxsDKGVQZgR2PNup1GpoFCv+tucUlA94DpBKIRl/1
4NEkjKGLqTuopH4e+g/23//N+we9UDouKquwDEFrMpVFGb8jIuq4jN5FDWV0ybiD
5Ba92F9iXGCWdKoxGDKdWRh4FpWS9Rqro6imhZ5NpuxKs4M9E3MAethCJtG+HkMV
kKywj3nFikZ3jURyh+KP2aBSz1lWuj4lqwvuk8LaOSA27roQn1AXgV+z1JaE24LN
9LeFE7DDLr3hZcQOYVNQY2JFh5cdavUWz85hLKXyWP5YvjGZfm5C3il7q4Bog+Ew
Tzkkp0XHPrpxyO8QHKwtHKhwMHxbmu1CtzcOhNGkIuTXGdRaJPwKdpn3LJOboZl7
pgr1gv0Yx6WsJTqTcA3IROHgta5WP+LinBeShG6slLDfdxpP35qeAgdaURsrvqT+
dBPfcNknmn6RQTKhO2i07LfPppLI62lLqVRk+jNtehVmVjJ9ulA9PXNs1Oy8t59+
AeSG8H2CcAwaR3IRfSTJfa8FSnMTqYnN1GU1apnPnobAiskpXbUs3pHbwtDXySqn
h3Mgcz9VbkebEqR05tq/LIRPmVjt7/nXZ2+MEXQSyGMOz+2p8IHSpj0Uj6NFfTgb
lYmhiUROd5mFR+pCp7ZiNOpK52nOIdPPG4OvvpjgGTCGHYFppAkwJClWAHNDGJwL
hMtDxUbAIYDoZrab7hAWH+p2D1+IrACevpxwR3A433ieA3ddh+S3yn3LCLIzf+ta
881kz2/cVgS4PwkEe2SUfxJjTHyhKyFUKhLwotkRWPXcGaUAdm80VdPcStIScGkh
jnZPGu2x9JwcELPaPfdjqFe4uZDnzEhHW8SdK8K+s/NO4OHj3CCRe6x0CdprFMin
XzzLIDoTwqIWroktKkhcH9OMOSdRSHN7e6yB7Lxhpn9osvJD5M3K0CV3wP6mBWfy
Lz1JfTQwCvjGSH0/PaUxcahHaA+hx16FverDRzqFIC1/OU30M1yhOHhsFByNsXxc
LDHlabSCNX+qyP6I2LLmU5R7XVH+DylXhaD5DKBAYiev2tH/283a9tv6S1+q1cjK
/yenFxM4xnBuC0qkMKmAHlXUo21pbKBYF/rZhC2JXPg9Z+6Gk2p7sI8Sm5aTeUPX
t5ppTZy8R5SkriVurXCximTOhJ6YV0TpoauidlU5knG2Zxxx1IodsVvNhUSi0Kh1
qTgqVoWuWHuryvY2Cy1PtC4KwPjt4p4+aByo51kl3MDvD2YQ+8qc2P6pjrkxJrrq
DAHCN1TjKDtAYEikRsFYKdreQxPe+2p8XK+WXG/rFSNZCR5xMMQru8VPQyJAlvGe
YcC04/FB4RjtQILX728iBgH9NW6PGixrCXSMBX3zXkCcl+/BKiyW3Gx+6LzFM6w1
D2Ae588cg7BljVJc2JJPvVXPhVirhCLw+7/j7VtTW66uQ72DgEtxvCx5cVmSYCWB
+n/Kt9VOmmY/PpNKVNaaNhz2VIE00/8FvaQwZ75c+iZU9x9tsH8MRsrl+YctHDsj
Gk4zLB/kfwcL/2NppvlicTnxQU7sbgjhCljSHd6KiBqu3B0clTM5eWW8IHRHE7Qf
L3B/9eXEKATo9jK/85b7Npep6nHQ2db26pEfHnbk6wZRLYDPeJ8i9UBeGmyJQVRh
dLaqDGm5Up2Zy5Im4AxxbuHpoG+JqXawhQYgAs/T0Ab1GoRrYZNWWjR/juiyq1Om
yK0HHwnzykHMfRmqbtX5+o7BQeiyD7xAwWPVlPNdi1lJAg5jrw1DdYxOIicYnMB1
6+adQt3L8kwUVJlkQzeK8KJsKuXCrjAg4+rSB7+SLlfQBMfDPWoWlxusMWnDwItn
hTA5myMt6dk/OnLiZO/56ZpCif3WBEXCTJ5hxzNdjGVOVQr4usbTOh+F2V/oIhZI
2P1k6tCwKNiCy4VlFWSbV2yYh4ZkCnZCbYJ0/eAKVY6qE3NtYSjuyXeEbhf7WPcF
xZcSq0sFkwtEC9Zhq2jSvBKLqP3f0sKoWDfeDKp36fM/nlm4BYjYP+0H2zde3ifE
w0wP5ryxYZlJTcacCdKkl66jOP+67eSY7PZQsYFuSDzvQ18VpoxDQSh+MoROFi4H
6GYnXTlZ7uT09MbbM/TNeQPzL/xCLXFVEnqvQKka5QmBDhJ04UZcm1eQtVIbIEPe
nq/l4srn+r1kVsYZMSxk6ayyaELM1B47F4Ttbi8co1h+FZmcrhdX9QQjlV3Ql/Aq
8zxYZzqS6MHQxjXvef9BvVXnRZVAwpDFsdL+Y2rEAJZZEyae+0uc2xD0BfcOCv+E
/V4LU3yO9ljATAU3WhQC6PNQ3WrvBApv1O3qz0tRFgo+wwVoZcAOB0HX7fGnxZ9E
dw9sbe9BLacAZVfOF2CFvwR2FFLvC40aO+QymHBAmka4CBM8LWI8WFSCe9jvLGKH
0AOjsFZUDi7RDpXoQFt6DPFNjEdhtasPb/YYIvV4p11QhRrvKWr9I/AgyXnKQdCw
FRUr/Obe67kGgZ6v0EjO86pHuYnxMORVb6Q1pmQ6VgNsKTqyUbH5L5xlqjdmoKve
QWPIk6rBLDLJHJRaLLUh7dbP25wXLDGuStbaK04Vk6w5oN2704/9sRQprN26ZJWd
omUHhZ2xtRPgXPEuDwU0JJ48uiVXtn8V3iLKMr+zHuAoyfJp3JvsRXMRUpisB1i1
+QTO8eUbsmZggbFfKox7pxkbrllxosLjyToFBV6/h9caBQSLYHetEFtRSkLckQv1
L0e/WfyJ+PgXjIJ4vVVldzbeKmdadejcgokNJZdtkm86E1toor3hS5LmycU7KgEn
L+qVoe25DMeqnFsgbcet6PVrEzj93TQ2znr2YtKV9eLSBLc3LfqgiDRGA5XSdsh3
m/9FYnIIDPcHbfiwDbKixNJW7kobQOYJNOrs/5b/M3OlpxbhuBH572etV4ALhneD
Do2Lt/uOVtYIHMwPT1O+9JjYXbTl2VCAI0NO7Sl7gD+pK2FIJ4Rj1egu4ZkouQUX
z+32awHhUCOvmM0WUEG7oBxcL8tk1NlIBHT4TiDL163v/m/411leS0VlvlO+FSAt
J7OprQBd//aMvdr/UwxPKTehR3Yg134yaw1dXBEzzAKmnhbg/Fr0o60tvOo+T2ca
h2YPm1T0ROzD6uMs0PDrxQ6sd+82CKDOE0XSRoDajbrN0YV3zxKfTodyPTOztZxa
aHZi4MvCbWkUwZ0ajP+rvaWKtczIPgK3Mo9UCu+mydBq3r3RzH+uYrn+n45f+Dq5
huTcfg+ogYzTIkKDseGhOCvOEz95WbHzLnLh8k/cTPAXnueb4GNx6/S3DwY+oKk8
sN+grO/5yWMUCBcO+1qrGPw5jXrxh8YboCYOci8v3RczXhl6jlwpGOst8Ng/0/Fj
9DXJSI4IYZLs4bkLrcPdHcJfmsmv7WmasHAgO+Y/ZarSK4QBoh5U52FyaRPf1Egx
K5vcbr/p9zyrQTuIsMmDr41B58FBKsY82exTSRd8uBJ3o0QgNIi4k94edio0qK64
U/MY9//uhO80AkiAcfvoZQ4e5EaB4i7iwf9S+de2WT5vczZO8e5UXMEBMey+aoGK
BSe5pNr8djPF4oNMJTeOc78T6xskH+JqDGnMnd1Oyof1YpcvIJkELaASnuS3Owgq
nHPcUx9LRJst8K4Z2L639XuiE11gu/HZvx9L7KUs/t6w7AztNZT6S4R5QJUHCiq7
A/x5BQNSuTckzOpaRqv1yX+Oh5SNds4Y/2iku25/ExVCQqSmzMz3xQZzti3WULAc
YIlz3TaJgb4F9pZMApsVfmKfesYIAqjzQfYHiCnQ9PAjdjl0M/XfG/Nvoj7hoExf
nr3d9P7MtaKq6vdtmgplE77W2QBdud+9HOfDWd+Irc+1jZZPxyJlYCxl1zfcFWe6
Ss/YJJ+y4n49mlVZIvo/0zqSJW3htSaHtWStppU8YHSH3yaavkZj3kRMBpdh17Hy
XNJMCOtHUdePHzVgZCnJXiCokQ4hjetQlvkCZL/vrCxxNQu92MxFxiQaK4kSwqhi
Tny8Xna3P84L1+mhGK21fu+YIdnWovAPxQR62U529ng4/6TDllDBhE7/+UKvQApj
5fOsXxDy3ASVJiHCjLOwjfH29P9dwAnvBSkpAlmA/Bnz1plX4W6StBgfSt4m2py2
89NBExaxSC+wIvJRfAoLXn8NHHeqxcgOZpY1RjIJPZs8gct4XcY2IQgdKQkaZbWh
nWyn/mwUhrmealm2/LDiZfkckD8tRCaLCzjPYLIX+rYENCrV5bESY5S2+3l7p/WA
LHKfL2vdx8wUl4Sp7lj/IcmPAlU1AZUEvfQuI6eKfzLK0Os/CRylq4MnyBj0S4qr
GkDeO1DYyfwU9VMK04eZKoATUz5m7GJh3YKeVnnpyyqj49QvZUUzwRL8H9kk+hUU
xiEn9yaSJl3vJyiBqmTc/kZnn/cptOe+g9ZZE46PKSM5KK1mXG5TBLIX/Dv9WJSR
OOdgkZJKpWaP0SnCI9qQ2K5cUsDFx0BSGXzDw3IhA5cmX6Zan6nj05AidRMm0hxx
8Xf0g1/cfYb1V2PABfhMag3S1F5vCH2XkJSlsLy4ZnafgfJW+i9Ii6erQYz6jIes
7BsyGwXQI6Vt15DHFKhJTVGaZKQj2YzycaFy/mqe/M6wei9kKsBbyWXxHnMRIqNU
MaxRDPWPktCKDr4Q5ekLg8Sk7i02zW5thTVEeDyWubkayOM7Twbu4byUw+QJsdnH
uf4wSsQb5fRFU6kV4A7zcTf76DPCBEFgBAMvODstSlhmL1ggB3t5jg18YPh3idoB
7txjTAEb0YHZ9ylCcTdaYEi/t3X96cnCqDJiAgiMq5KTs/onfJGLM8E1Aoc9ySfu
gEu5biS5jQvdpi/TCaq7lcBSbZIN7VjvhiMtuLWT7inRFw/MEDaTrDjev4MvsuiJ
Bz3OQTQIaXJiJmNoD5XG9jNl2sjto0VwmnptDuzODG+rjokUMRZcW28/w1jXMmg8
Xhhs5UpZ4tE545ODMTISoIcleE/4xmwM+TaakgQvSiHcWUi/d1m8jo89M+gbcPgA
uuC8jzV1qd25BABd5ZMCQaNp5zHlk/k1sH4Hi4zVy90uyD2bQYx/u8YMC/4EF1lB
a+ynbpZVPC5KwmPSZUq6JsmwHOGclmphpeAhqBa0bP/WQrcPzlw1099CN8il6KoJ
8YJfrAn9ajDWE7OJKz6tX3dzbzheF7k4Aond1Tc0Uvj3UsZAt2W269TjlpTg5y2c
xzMgfzRKArMaBhanq0DW10k+89u7m369OjBTZEwJjVIxVXS8nYas3P/DBjjnKvJq
FeLrxN7BjzW83Yx/kij1VFHlg3ypHl87LwE4pvOKeLEgvdkrDAktlQU3xp4+9dos
kVLN1Ccbs882vbwCjcGgRPEyumv19ATC4/YU9ThGuJajdpsUNyxswzrrR1eSNjdD
7ONWStSLVAnS7bsLgfc0UApfbHhb2Wsqe4cJ7EhnPyiKutTJ7p11J1IaXmjHndcU
AArtpfvYwDlbtevwuuVh3dtpfEomAY5GZgvEeDVT5rshQ4OMq4jv7OgelcHkSD46
mjEPugMCnHvzDGBHsRrhMCAG4Fwe13KSaM+cFAwRz27hS9I8ULVerKGBxoNAJQR2
+avvdO2f6EKiWACa58D9Bvj3LLdu0qX/6BZ+m9v9lm8ZuU9lfqflx1eUxgWZMjXO
WChbxdqiMqCTeyDuxdK56mflEh/2V+V0vMWcfBbp3x3tpDTNEZJyozrbmMUECTcz
GG7BchT2zRGpWSgH0kCL7tEVRoMJ2apbeYvQ6INbtxVreHPUQ0rRr9meczk+N7hI
DPQRHjGZC2+tTGVx6LOIjKa2pJ2q56jZjZT9oYIXvORZf5Ai1sf4e7VS2aWdoEoK
/iMzNDEhQP/9xj6MmblBb44YzvhPCUrbyttyuxO/J1WTF3vqaUJzZyu4uTwldS+k
vICsWmVNL2pBr1Z7GItmpV2dAw0xHii9lMEGsDRYhgmRvWH7XAPfSTRhd1KoPzFU
AykKLV6Lc7noVsW3Qpwx5ZpI+yShdrSLz+baXZ1RicUGb4WmJ17T1CKWIOAzSJCB
n98O59gIWntvLU0gtwrk+obbs8IEcMTcJDoil9Gvcj8u8a5xO+hkI9yoxYCkbFp/
Tob2b9ww8kcU2zV4hYI8P31myvUB6WFqf7887AEsi50b+l3QBqHYM4bBXtwSZSag
dmYEbboJZLxAugOvur/EGL/2xzfGAs+8udT9ohNZ3Q7RSVxwGTdcRWEprDQx7lkT
VF48QWjbiudQBkjud/+602ip/Ww5Y2xIxL9nEsiFL3f1+3YPIohJ44N1hgtW2pIv
x112cMfqsrwX/ytlbbY41q97Ly5m/Uy84plwTe8FlCblMKYBDww7uUUazIqzSump
3aUJBrpvEKtwhFj7H1E58qtOHNvLWuULB04XgReurSybtE7tmcqXl4G4EMjBq/cY
pyGlGdAJi4qUQZ06R2V3xUCs0wsa+IjkSg7LjWb5u3kF3b/RyxidTz6sP7feQTag
gWxTixr0eeBB+jRrwelt1F4vd+N/BiaLLtXwqjhFbP3LPC8yOoBMtBDKfPeMM9VB
lKvIit7xPV0oSwsg1t2ejFSF7FKDHSrlCzq+Rmx3YlKwIm2IwoC97rsIPFvgUwwp
kvH2CQDvFpoFqIof5oRYTvlYC0OFni/vxDGQdcEANb521iWt957uj7hc9L9/mFSs
lwlQwbmfo91cK/6jd79gDRu6EplpYgL9OB+wDehqWEnRE3jCYyYaENvRS41GMCdk
mWye0Faa4/wYD+Mvz55F3QtGD8m2bVxdqM0Ew4pzVb0wO9ev6H7gPuhbTqiFVHY2
WKzP27etNhfgjB0lUOHsj0vkszpmCNwvitfO9cYIXORLjpDT+YzPlZY7OsnoVuvU
LxWbBtg36vKAhSRhcQb9itLhyBq5SJ+PAF5JjVR48iH39AZkjEKgpYVlnmWfE1BB
IHZkPU1r2cUDUuqeY3iZshxBiifkFdYM/84Pt6W3spIYAAe0l5Lpv17uaQaNFOeV
b7P1p3wQIVCfMEzq/XKUD+hbK5dpg1czHlPdk/prCDmmhHT5P25B8X0tzH/A/+R5
HMH27sGmpL+cHnAf1AGbHces3cIrRx4jh++QL5dSJQ/Lfrn9BALSRPer15F30x+M
w83PhVXx+j1GcXLg5Cymnyy3dX7f7Cit4oFb2CbyEJAUOr6AJi/Q4H7zQ/b/brew
hIDTi+03d/FLvT2o660rKGFUzb83ZvAq/hCogQQjZ+xHSusgxi1dTyFZ00R3U+QV
732VygqtMAzt+ioFxH9A5mi7lJIR8ZW1TI6lwDksF1egE2wsOj2krGsWdzJNiGfM
tlYYffgUkaHfhwk3XCWs+0SRBjxl+3RZyDNi0owJlZsjVgR1HLq8QEChRYkbjM8n
1lzngRwZ8YKBVTRCX/NFkLoD5kUyA6AFN1R24FjWzEbOKxxTu5sQhlNN4GiqcXBs
7fTeVGDCNRGK23VoxvY0CfwX9ivZ3SW9q0uSj0kTyQpGSWr449q3XevfM1tLN/kN
NmBrBOzwlShfZcB/6hBlXT2J3kzPDUxW5omBPu9BQLKd7T7Zx0DTLszRAWwlibZj
xDDm4hTEXhvQC2TF1dtsjP8rO05SsJyqvP+DE8xl9D0Cnl4fdJ1BrbcI0WCd67uH
1OnA3T27BmEL1RUWZUXEHCc4IQRDZ3rDPYpWGlbsjiPM2sSj/7vaJj6Vh3G0DTDT
txZw5vt4YYGz8u3k9yS7pp7fDI06h4HzX6sTXHXlSi4b2NubfoSjdyfCM8ZbgUw3
924hNh3Y+J1bNEPSC30Dd9BgytenFL5Y5HsZMtDK+1PD7UQW0JhG/ge7TpAJmJZY
nAutGO9dwnAZQrWC3uj9f2461gtP1yvX7WDWqLt0tg7hwk3Wc9ddE+pkLSFVVKHT
vHv5Zu4NhblvWxZL8YBLx8bEhRoMWG+6ydrLpMHZhGfPPLEXrSa6NJWJa0fDt7/i
JPfOko2QVDZL7chiO6ExRQXRGQNyTqWI3GoqjZT2ODwv4+kkb6B1G3BI1NaehMBG
2LnjIt4B/pLt0rWkZjPhVNLKeOt6MnloO6KR5PA4Lp1KDkTde7HKvSVFleifKbcw
b4jfU3zzBKy2TIsBq/XMZEON39ohc389T/6ILj1MnXp/2ejBXrAIf2rdULB4DnQp
Qj3HIMqOgxPRQGECUchujPQ8pIsJy5m32p537pqKIoUUs5wv82PqVepoBZygCpN5
lnxKJOyN0jDmwJkcho36BsBqJ1SpH3/8q+btpazuhZzRjBAsKYnNQ/1rIXEhhj5S
EfZMIW/xaquMFDqBF38dDOpfW0uWAGcMzlR+pxbs693f/En1aPTby+UAwbRrlJyz
FPa7hmy6qbrd2FfWRUpdfV+idLjjwlXjdH2j+4xh5Cd/zrApNFa24OlGrAU+tAZW
OFsV9joV2/MZD9JnGsfSOq8Gn1WZulOfvyigk9eig0q7DiNOSjxSLXg8MG8X6ez4
uj0A7WPhkJdmqFhSokyXyNlipkc7OmWf7+BmZvLdhXGFN90SnxaHOWhTJyjgTlFm
lpedXyMU9yhxC7zs1C+xxoL6uL4k2GmgmPfSrwfCHdz2UU4H6nyoIsVFDerIowxq
pDwgGpBb3yO73OEgq510QGMTKearBnkFuDySUSXpzFzO2SY/goh6QK9gFTGnrU6i
6QNx2yUtfb2DP4yhKHD+LROD6uxEStvvnnA6mreKvL05K3FzUPodVmZo+BYYIplq
Fj2dD+oRuMkSZx+p9dujdL/wUYBWwkehsSFU3xYRTsvRsWa3AqhqU3mXxzJ0Cqbs
rn4EVUKue7UNnYOlGx+Hi6/ozlogcdONzMn7VgSnt/1Mhdj0zJYT7XQp1ZSyxwa8
+Uw6pY59zfkbgpn6KLYrShZwYffsaJhaLoTSKli+pWUr9vaVhAT6NniTbDWgkuYK
JLFaUwR9atT//tj2s0Vu8yOiEcD6r7wim5AUU/RWn82oaabsdbUw4FKLnJ+R9T7t
1AKpa3rU5tPkLlYMGjaLZfgROi6jNMfreg/IXUnsPwlOyp5Ku5DI8VUUoJkYh3b6
fkOIybEtWYVP5L9VE0ezd7OpXujLpe9Xu8ZRsTZVFqfSVWUV/emRFTvL9osj7Slc
XkPBLvEI/kynz2kG5hyOY/NzAHWMqFcVaSikAjaovMofwxmCjbXBiWBT4KtEEANv
HH6+rk75Z194lIECx4op6CCsp4isPKYPbgSMWMDBpgUpiULK655eR9hD1AClEc4R
4lBgBuAJPlYva6GBu2VqBauh73haSAv+OF7ugUKQJgeOtQIH97O1cj7Izxdrw7va
Fq1P8wsLz4uQTabYd2Y4w4oMFGFXXeu1IV9+hi3xsg78LKoe+No8oDT4hKQSywho
ng+HfDzWaH99b/+tRGtzCa+wKE3Rrc1JgEMJVYkCdbw4+LgZw/xofahJEyYHW8X4
5zemKUF+pPCTHwI/NaP+vxr0vlGlRhMOq+xuP4PR1XtsoxX2zi2xq9VPfTvDLD+j
GwIFUnlRj5xzZa+W1yJsvXA0EfZewN1owEc6j6+zcLylhimyQGZATzbaeJ33Ozu2
vcPN6mf1Vim0ULQ15Zp0Nj7WGVMellSeO9Hvpe+UsfS5qBbxMYlEcSnJlHEv7pRD
zj2f6LD12jHqb8a+Xhv1Otwvdp1GV/597XKKLcuuPZnHa6DpUncqqawR1xeyF1X9
vnyeLMF5BOn0ssCvAtAD7RjUWhGf5HkKl2XOPD0QeIMMv7kbU3PlZI53oKetT3Le
Hv3azxFc1uGgR7pZzi8FJrvm8yatAgVjNKxiXeS4RGrQR59KyfT6h3zVC54HJhFg
lU70ZVKNTJaoujbh3YWIPJMyyE9Z25hYrBM3AQkNwlkiz0y11hzsmXvwJpUbhr7+
GbnB4QpA5NLKLcoUxeDELAaIYVHwwhgOHG0Boa3uYGYfgM9gNdCrF/mTgP3LE5Lc
tQPLs0Yv7iWBSE2OG4escdEIpIahQHwy4iZbDRe8BEaNncBO84Rlj4VTnqdchE//
9TQprmQ/MmvV/rKhnGTeqzJpbAQk1GGXMHAs13jKLNOWfFevgfLZfo/yKXUwbj+N
2el8l0bDu5f5sy1EHQoE4rGDeJnkuMpkt8W6pzYjGG+t3eGZvfZ0NVee7iPC6yQH
nMzJUjPuK/Gr1KMNvrKJTBzvcmVhNGLjIR4Va9gCA3LM+uMrIbFiTVq9NxFPkIRd
ArLkh6CGScv+hBGt2NONrcuMi6LKAfnxZolLYQFMZgh8Um5JE/cwK1jq1nWLCsM7
F+Z8wrmhoEEPZZdi1Y1PyIK6fmBm/I5v0gIVN5hFjUFmKb8ZNVKfAbRpBB4qSC/o
plfEcMzlVXUU//pg9w7TN1NRGGI9LEW5I5dVeVeYonfdKcUg6Dy6w8kvxaOCYQ04
YQwB76eRowJoN4GuOB29BGuSAqQp/xL7sFzzYm/8opBRwNAbQaY88CILZtIKbRvH
bJipqUGqt6g0A9GIWHJTgEm1ISghXOPh70LJyqrgxe/Vk61/ZiEhPUcDxlFG6O/S
KwW8B7kyPdf6aFP890C8QpNaVyfPLmGwPYv1Z91ibV5uD+OGjDihcdt30XvcmNZV
taCXMybGrzaPN3axHt7KSWyGjkHXvVaKSl96ufcU+S/isaucyxZKtCf41sZK3qv2
CEADJJ+H7oy+kgwROFV2MyV4/XaAzc47jJpppZdVhlyCyAVMtYSJL4QOUoH69Ovu
uAr558TXIuUZrxuBchq8UHc+8aSX6gy3Y4CDFQZTZCO+nXOe95KhzJYSHH/1dLkG
k67kJXro/F4FxGkADu+476ToM44ieybRjBEsueAvI002EXjz/FtM6qNPWbRoBRt4
EmGZdIHS2sAX6oaatD5NmwwgnlbwJNjA9sNlRZYTMrioy88q7NzxV4iA0LomJYi2
QVljWqFLHkaJ+xPwflT8lACPocth2lRV8wlj/fyb5IMCg7E2fP9KispXPHuamTfj
QFAwBZFvsvCJ/icoWFHVQ9/BZk744B/fvNMg0f2hH34Y2A+NxcpOhSv8OxLX7Rr2
cCnT3GQ6pPoRciEkr781ALKRqUX+ktlvrx6DOeiCo//x2mxotL7zkJaAOY3yFTNR
X8XWCQo8O4DtnU/oAFcbxbQsslCcfdVbOkpfoQhlCy2NoX6I0cuul36h78U0rYK/
PRkQkoo/J5F5xWXRya0ftzz07xpXQMMldbvUHooSiZ4PObkZ1+ktfAu9RsHmSm3B
AvVFrQzs9RdLjNpSGh/cfXCL0zH/vNYdTUzLbkNDTPg86Nevq77gt2jRjqSadVcH
DcsFLwsdfNQE42mFBbA7eObwdhs+n8tjYenUFNHwNznB2/nzUKuGSHhvMU/ApdU7
N/XgqGSk0jqqTjyFPCeijCFR0hLIQ53b04pkg81UhIZsQCFlLK83XAAgGFiZurkH
ip8TMJw4aB05yXVYPm9LdtA4OwdJzpL9/7rq+ZrIF6jmq6u+jjb/I4ucC4a8Xylz
df+oy8y3IEAqH4CmffSk9cAHY05qwVo2LmlfFVQIWX9lDA7fdNKMRjHXbxR82Aff
tbk1xezaGN8WIPVbZk7RBxFdZb2Wu0KnjOfyERQ4eQd6GwzDD33se2vEzB+042ax
PlMdd/7Yf4HAkO3NPYCvsq4QYMIkHworT2kZjae3FPSLMsHAaXn+kdrrqcCRRtlT
7QgsUgRIAahZNwBCqjUWp3puFulChaQHUGIDoJt1RGDe6s8g/a4U9El4+4qmrAJR
fzCu2xQ4R5cs2wNmZzyjBggHnHjvIR5rnz/wsKJ2iWj0P+hqD4qPMweUS8E4308M
Vb4LyRZtjvQ18co9800vIXpMh83RnlKBtUuiFUHuIpMybkAalHde4m2C2KiIMW1K
9ZUVdaBL9xYyt7UA8lEiksut7k/XauS48sl/PJsONCl9mivViEDkoM1/cnYHFSGw
SXajnsbLzL7Bn9+bEQcrGeHxmEPpWqAJXcg+dLiXUeXhXppuyzvEp7As847GlTu4
8Jc+gTn9V8BD0Gy2znl/+HW//HKxRfCVe5SDBGTOzlyhi1DHAvCdsS0zMscoi6tu
/HMEl+MxzH1K6yYaFthE5lT8WLSAXU+iKXHKqmBtHRQ3Pw7tCrNA/aqVSyp0qDlx
ln0J2F1kdHsmjXHN8tX2rpJGplQxBtyX4pDU3fXiTflr9tJvOLORHeXkdGRMu9xs
s4SU781w957bz8qFdOr0pbO0E5ZHTEuD1QrIPY/2tjMuUWCR1iii1u7Q5AO6hlsT
TNFqCskxn04RahNJUSkhtCN8Ve7dkntn2HVqkaL2jGTDRdKFKphLKNLoEBtcw+M/
owquBdsxCxRiDpals9q1fAlF2iCuumm8uGnBmdnHBSMUm9LKFY3RsfweQCfQquPV
Tn7RpiN9wRO/KbiKcd46sFEjLpeQJZZyG6VY/VFoy2x2oIsRY0tUzjnlCOM+G4VX
Q/FzcLz88TjjPzZZiN17J0RQpKGlWxYMa6VJ7nLsXxW5ylu6aonga3ciUsciVxzc
K1VA9NBd9XpFEW49dy4PdDgnzEr60YLU3aNAoaPqi1m2NeqWb9jhFApd+yQU++mT
toiO4N6h5D8WaysbHprQqVuNo28yyHAWrHL0E4uQHG8S0D15M+FZKpO0BBSL/vRT
+IDdEpcXYgcy+zFwHKgkP6pxyl7DTcjvOTfi9hyezoh32KpB2sGvnsi8gBDXkzNV
DNvabpEeshWu17L5zT1vkUx6GcNK85f3KyeLW02t1dIk5FVRvA6AWmxDjZIshB0S
2HxNwhAO+51lNT2pgcKwftQSuNLwKPjEpBZeapgllZ6BzJD/coSJBQf5GE9UdISg
V/QCGO9HKkPnzhcruTBu2obAWtMFDxRbg1pvUpX1sBWvvq6BZjj5gK7gy6IJiD1E
sVR29y7byTqcZNeufYHRCqsH/ly0fiAWIl3NQjr66fCCrnqkdPYstYlsg2gShEEK
eFBu47+v/tVflWJ13JjCUn18ETUrjs5eITsk/bWd1Si90n3mY7DEP/6bugBeOeYd
pmKkMDiN/e1FN/MKTem1VKjtt+HNCZaR58cx9D24V5Io2ca8zOMvouLKrBxr6Qvx
xqmbaxFteHEcLH7W/4GXqG3GS5j9d4IL29mqcaKlNW02l3MQI/mMnEXAEUT/wIhP
7VY7hwJTXysErZdEDWmZxDSvno9AFWbC1iDYOtzNYneiStciAsVboR/9hutG/ie1
AMrZ1L+R/00/sy19fAwK0MlDhNeAZX4+6kF8ck1mOeD02zVz9dbECaf4x6J/i3bc
7r5YdYO/0y3zPECmwVRC9zUi7VTLk27ccMImhfW9BAa7t6Z749IaoewANYl96EDw
Xm9ML7M8hiDotoYISDMt279gIQghoDP9s1xvnf5G0u6O91k9LnYjVdLaQfOVcM91
AMz7pkhzyeul6OmioQ+9UTyDGJW3557U2Rkom1zE8KrGBzAcJMm9F4pHdgfZo9tb
Z3uBuHgx8vbdMqG/CMr4fuLnk8y/r5+BQzbz6YwWBF3A+gLmbEFOoBdvHlgCeh1b
j1ZOe/pJPyAfSqObzDw0Yy7gqeSyIXGUUk5GdfQe0JZpe6FYW2sew0h2vz0Zly5J
uz6fb9v45Ye42WFsxBap+fMw/IqTuf/MwzmzQ/6GeTYHwCyNss6wHcxipHukprHv
XxovUzkz3+F6Up75XfygT/f715UeOvFF0wjxWhWGwVXk7T0glRptgDbI/xvrn8Zd
YOgUF/Fhzn1hIzCcTc9f3kMW6mRxHreAJ3RmUtqvmvJET8JNDAfu5Fsxam8UHrE5
L4PbwdsFEeDjItQLm9eSvcHG/M9QQt3YgyqhqmxZtTllAlSnEHN8DJrIJbtsHg2x
MlTvA+IMXU6ANnaK0mtUbPwZsZkQWj0hM+6H+eYAinXR0NWEyWcjP4b3V9cHDVFk
o7e6NHMvcgACMcVDwMm5S/C2WF9Sd5nfV40gwalZ9iV+fSN+3pfQooT3k9WuUHss
vVYpAI9NTwocb7W0d7T/KTJhOQ+NAfscJXuTzvzKXXqPlFoqRNF02qcFcqjtyK89
THd7NcMkmyZ9uAzssyxWOqkhMRB4XPYnvfy4toaJpaBiF1WRSdoPHFdC3sVUvmYP
NNoH6K+EIpBv5WTAJ0EK+mgeJfwlfZSqlq/GVSO3OG1irpIHL2J1EQfXWela/wJ2
cewsdROLQ73Y0x/lUJSsqKBBcLFWTeMxBNTVxI9imI3qSvVEjUAnjAS4UdmYPtdc
gBaXBZ2xuiUD3UqjczDR87xpiWFVKsPtHLHxdwBX27IOra6i+XVFP2qYlErrwp5w
uAq2GescmwsCfs1eNXuLv5sXP0USSVWc0HWs/WFxf2H3nsWadP9N7/tzTrZ9gS13
FJzOTr0fwce1x7sKoAiExZUYOcHGDvIv8ofNz0PGOc2y2wheeFWVMVlnCY9iokkH
MzFbr4nWqWWWYOOLbEEKKX/aR0ujvqTWOamb4kQ3I29E1OV4jAFjw1Nhfsyu6VfG
IwC6miEpcE3zs/m6L93/8bjJIe7DKbVVrLfYEPFJ+p1jt1pmX+ipTEYIcoZbv+06
VZsCTciX56wWwIh7Sh+8A5aQhiOqOyUxF/0rG2wtz0NuAEraKVVhcQV1jRsP+72s
NvOvYebqKOLQbpSM/qk6cIdW7kr/wzOOuO/fcpcAmv5PeOEGuBM6p16Z1XDjiqew
RRJsk3bjC+R60wmV7oV7ujsd4tNa+1+I5KdIjIpeq5ZkXMVJOmanB/E/Dk0eoyOo
eJha3GbXuaPsLYscnacjJOf8GmHq/Q7jw2D8+HKds2UlP+kbsS2jETXnjvO02Wyj
2ymHV/+BcZBXKYr3/E/isdwU11+qmSUJndZa8j3MuWsBTvxqm57cwQsI+6fk91xA
PYfe+UMd4oWFvVmszGr+ddKwdYlBUiLw/unRO2d5V5xSZzNxlk6uLTu/sDIw7tan
nMWUwh2f8vtF30TrNT5D0dbgsYVFt83R2ulOGjfqjE/YA9c+Kkhxo1NV0UgJ0d6r
1T+LPgWMIBZKgp9DGrxZEd9obRp1FpZIWj63wWH3FIIsW6gez3Db4QVs302AK/T/
5qLxeBxsWyNFwpW+nUc/5q0aQTV4qsanqa6IP4DPe+QjC3xItJ57jenNJMmbzB32
pr2EHxI0pK2Z1uOLehCe143vjg9kjQ5btr4GGpCkJnddhMpAr7RWmeP4i3eGdnd+
A+wGirw5SaNr367j1IJfoxr/abru9NsM8S78dnKk7aeHyNRVn088Sqo5U4QT9ISi
+QMF75GpkF9o0a/On6l7ws9lWvNACHVIIrHJxmlHkVr472VqLjeSuZI2CgWppDOs
5YBmSjv7BbU3EIk24+p6tcPurDXGGAt8N6EL9lkwAAm4udK2ujdcWZa7di3mqRrV
1Mb5m3ueXrxvrbtGUvHC2479TW2E2uw/7eBqHU6FSXlFm890VZwF9YbrgnNj+EnW
/WrbYHtPIYSIwjj30+476tWOZX526BAKCloUFvn6QeacNIOCFf7eEYGo6MyhrQ3K
OVfrOm8j5f565ItS08/GXvyFhK7l7egv2S0VdQXkj9q9XkKIdHgnGG6cn86Kiz8N
dUn8uVBHh08JxQQ6d9EYdMqudHV49Em0aXObrGYDAQTcaIfCYLY32OR5yNXgKdyk
UQN1/daPTFW6u0KVKTNd+zyR8p3pLTkP04GflATHGInNh9SVOgWPmNiPy+ilVrKt
Alc4pnA8NXc/KYNzk8nb2XFIUNgKbhRX8l5F5QkUKPuNIlVEmgM6udHoOAfYITRc
nrSeeraD8vyhPZIH0oS0gy3Wj0X3sDkJPvCUeD90vYAxvjQwQMUXJqnVbq+F5uRn
jjGxyTU6gJK/+A2njxfAopP2GxamZ4allsh3SIhWrmkOXH4+2TD2uQ4YhSl1C58a
ziDeV0RaK6Jd3roVbtcDpABvpKzqSVC1NdJujTenCRK9D298c7ZR+HNSC0ycdeyy
LS7XneHQ4DgE4WguRFvOlp1Gz+POktXAZA9Yx3yhfDf597/T4lcXtKvKFX+pMGe6
1VRBBZ0vAO63pv6Lzx5LiIlkk0TLuDiDp1LUlHevq/53QQSqGb/XVM4HiwObssCh
R0Sq2044TgeBbz34PYTgsGSmIbOLzC46hLA89KpaS2eVDeaA//uYurKstK/AkuRw
pXbDfLE88V1YzkMxQC4j6qWrqKoK1MS5wqLd+XH2VlAfztEdi7VSfamDTtHvM2RK
xn1sw+5nOL0q9JnlAqYD9EVIX+Vilf0dHdtbljGmZlLq4FzSZwp8ren2EsvE+SAR
0pWeJKmQjaFa4Q/KjUSuKz5g8MwOLx4jF6gYmyR+tVuL1cA73rpUWwNern+FaIz3
Tts/vFzJ+EbuCO5mIPKiz7RXn7boC3V/IMktLTxygT7Xi+w12GqH8ncSydzayAGL
VBTPVIgVDBmB1Vhk7eTqF+bkiL1bTrZbQVt2ldMDvchu2BmCaAx6FSh4R8ofcGxI
dBYaBSHPp99+8P5PboHFJ+wWKbSWCZjLxXI0//8l3NxKHwEjZc1KVH+WBxYIGvmS
wj0BuUxNXmLdE77UO9VNewqA8og0+j/7/7gKb/dGih5osEnVqvA/ySUIa35oB11G
8SSLy9IkMFbtT7O4cgUEe/042PVBm2G1pdHJTFmKLCW/nks/nG/BTVX6aWI0HLQO
SrLQh3GLas8JpRzn9RhNmAfCPG8cS9Yyr+s6xORXXz1yu5xBUuar6Zd3uwuadIRW
p9Rq5XC8UPMstTl6gFd3gPUqt4g3W7x8KBV2cWhk4Jgn1s7/mwYoTUbDeubDaM5r
w8AobnKxRXWJmAxlWrn9S7VNlfH4FJmW3HWXoiZAV9mTFQQQ/q8Ze9iKlNP+7MPo
n/DumrIQn1x8/DVL5+VMTf7q6Ayqo8/PocIbGCF75o8xWma1lHkbchj68yhD2y95
BomZAuT9hraXEki+3kx6zB8tglaODCAiWN0/dQlad7jHJT8vjMwR6nUFHwIhGBrd
box+KJvqFYFBtW5rOnZF58VD4JPFp5eGt4LTAX9o7fpN80KcLOvy+Pt2kW1Jqxop
JmYEw85D6D2rfV6ReYwM51rLACJ4P1OV3Lm/A+BOaxr9zm5hTr57nhIn6sbb2uA6
4r72v1Ime4flglCLxbRqG63MXSgQwvNTHw+vOqVppc7hOgWjy56he2JZVXN5SeWw
XGzVBjaReFWgpfpzjrDybn/bLPuq9c6cGXEKJ5uVVVQLCdu3yHaBKpwS+I0dE3Y6
GK2JmzAl5Xu4nyEPjjpeoRJ0oY4wVHaXCes7jBjkyLbZZvtnchcvuUASe2aRqpkm
WWZ1GN7kHWRFf7aGIKGzIPgIiRo6oYZJOD5DIKwLz9DEc3oMLeAX6Na5v24hUvRm
VoWCG5GzXmlS3sf5m2c6vszlcqg35RxealGLAv2M8E9qldlCfLEZzvFR01l8NJSA
QqIX+OWAWsqCqWIjgG5ie0XWrFHmsn4ClXVPbzPObqTRVNEv0hBYjX/KNPamhHO8
5EyrGSII1NCsW5k+7QVSDP2JOLPtkq1fp+5pViJokV9AOxXLbiY+iK8vIrPFidaD
LLOxtOvYwn1t0NKk1FBWiUWYAL9EnzR2X7XSKxsSNof1o8YGPagL4WXNZLKV1kLz
YW5TouAIdfroU2UNRQQAaydug0FySjyRx7I8uZmObHASLdOjt6hR36i26DaaTGgY
/6QghnjDlAWOopE+P7RKbh++9wEBmaXKO0o6kZ48WLG4Kgh8TtzHSXTha5oC7S5X
Wdho4yUVTe63ZmNfaClknR3F940aLiNcf9ELZW+P8a3QlQjwKL5EOtCxtDqmj3v8
3SgdPWEAECb/79iI2iK1kIr2vuksGErkzop4lnoAAiyipw5KCQ3jf+wjHtfYUdhy
izqGw9HlQO6Lm++7U671YNYciXJ4p4qTriPZiF7ayeBC1+WyYWWuGk/AbHb3j/jt
NHXxSbAveCbjPcgD87jqqzFfmrGxJ+FgaND/Q7MYSf26gDmrxC0C2bIXoGVGneul
CnrVJUxz6AqscnjW2uFemuJQ2qfvYjUdVEtqlwLt9GDUuzR89p30f/z4jHL29Lnw
AX2TcXH0dw3KYZqEGJmi1JrUc7hvsuBdU/S3BhZS68pac0XEDH0dXFJGvW31CpDO
gy8zZgY0R3rWsRtXL77OGZUssLh2SuvAW6jev9ifmPlAoQIxiqJjkvdp8ynw0ITk
/MetPp3jLdu/+V/OnlYhmTrEklH6e2IifejGBumPOczEP+YlokfY30FdgWUO6lMx
s98AJAKGafn3nlzNBLxV6nYO+gmX6+X9Kq8L7auwjYtYhDCKoiC67KDS+WIJUIqs
Ya7sLvq2prfmJcr8bPtitLh0KYlV/NTXT3NYphOq5c1ffIYJBkqHm0sbcgEZp68W
HMdZ7BaVrC9SoIXMKSNZjlZc5Z/0SEgQcQYLjLx2JXAkfIHzkgI8AuVtkYxZK7Jx
1JgwkboFaBST+6etzq7d1pmly2diRqPlDPC5hoyx79McuScTn1nqPZFwMdVLeS3a
QkLcRfjLBFgxdF9a7bjp+e11a5Tm7lgaFGSXoaF7K6t+0XGeHzsORn6THDhI8WvI
BEC4ygwCBFn9MAL1AcZ1avh13LLzYFkJONjizDH2Xx7v/y4kxFXwVkuaWM3R743b
l6KwhnaPnmm4kNzlDoJ8zkg/4PmL0yGFDGn6VXwSLH1StF2nS/G4Nu9UpdFAq4c3
AMe0Jp7wQK4rBcOgbfRXnKyg3SLG9xk5jNTcTn43z37kX4iUXR+XTAyVSenOzAWF
iSWDDk3i7N3B5ZYo8mvsYtIiPi84g0QT3m8KL59gWCiuNH938KRBOgbSQyqvfswt
mAEYCFj4Oj+bCSi/K8matUMAFM/es5gra3LwY7pER7r6czhThzUlVqt7sjlegnZm
X++DiUREq145dAFFodOyyv1EO3sKkH30d5x0wSPMWDlfjSzCEbDo0genVPEST12d
IJ9gGTyYsIVhP6rMI0g+VmHJHUBU1s24rtQekWj9BddG0EygVmbzGyyK4td4e6Ta
4JaG3RCZoPUJXrU/G7Ky6Rc4IImSGCGKwIaxqbDx3CiCJTP/b0AXQE+IJqBFPs0B
WwNpXNwP8Kk0KuYzHighAJUUZalon9oKgnyTPSnQ4Zr4o98HeIZo2UfKV/qTDYcs
eL2RJSLRzbUZYSNQ4MXopzb0jRBdnFnCPzDJEYhW8oLr++ZxolnaRIe+zZu1teRu
UXP93kfX8fCh5Xmkp8yEiMHIcd1Z/YwKMuwK5NmUXk/hHNOXdOCpVu9LYVQN13VA
5gWoBfcrIMNOtCU6aQ/wtH+ZLyaWQhO5o37r5YH1690gPhmT1e2Zm4WHzr9Abk+1
IZ+/SCmLUP1hZgp6FN5qJ1dMayEFa54P9CmFwlu0Ev87jLbXhBF0abVC8SRJHdw9
/R5dej31G45RPV+xnXDM2ajiTuLAPKw49E9DwvBOwhW8h9yioN1AAWIq0gmiSel8
EWolsVtxFCZDofhrBBvPdF7yYzratCtVoM9ftJGH40Yf3LN+6lcX0fk6oFZCiMp+
b2MqYjXaqlGwC+2VG4Is9rhxhfLrbYO6fSbqQ4dCqgC1pXNE0GG8Eik9OlgMak7B
RusV00j5K60/7bdFSRE4jDXPZ35/iZidyZNm9vTxbrORI3cy5DGbH0dxRB24jrnw
bZmE9JVPYx6ZFmw1/iB7CseeTztMed3UU4jnc3m+AOmOzjfEsYLxCgNzaiscCa/J
BJizwSDdiMZm6Hp1hY7Ycp7W4eI/Lg3Q0ZD/mXH+9qnI/YXuNBaSrocwFztC7oDw
hkuk8L8I+Mx1TnOX9HpWJdD7q6m2DU5w0wBaa/7johUmJu8cFT7qkXqrYQxCOhbS
2nwpkUe6tEa+ECSiXR4aS3YeZqDJc2kBg920FHAAIaHhRup+Zw4GufJxucCRWTVY
wi8yd7b/eKSgc+G3LdB3dJbGYCqF490UeigHa4eWIqLQhqTStPQhTtji1/VOD/t0
7vlOug9OZICamUqMM1JyIO/bJh4DBEo12uPEHQuAD6JNRL3M0YZR/vJKFRcQsg9v
FvPBWxYBkzjAT42O3W8d+3e/v/uAT9XmH3q4KvM0NBgi+GAzeYbfA4t/3X7qPk7E
LWAyUqPafboKiZGHPSf1owJqHvqiHl2AdPARMuLNAhcdf6+jtyPdeO/vzlsgtnbh
wbS0c3ctZ8O+yY7RoYCU38A5iHLzwGhzqcLCyy5jAkq6OssZ9N3jiu6SsedsFUtJ
qLrqHn9AhX33CJfwRV72C2HXytHACgeBlC6X1MQW4RcFHDHeVMgu9MlAIw6GZxTB
0l28djTj3kRrMhnEAn75UWeJJFfpYQlfscPKYul160po+4sKROqdyfWcJi+8Vsj+
GIOvfszTelhBI+AE4mLp6/DE3KFyYCfUASQnnwb9yp1QxK3ShC/tgm1nqsmUifQj
aBgQWea7XDAmMYerfOR/4OM66FBq5Lic8KxUgLnHzt71QyhTANJ3MYIM6ACF5RX2
FMg2ot0a67Qsy7V95tXynkGAAoNoZB+568h/cBM+2yOFpwK7eqz/wVXUcK4jMpN6
STRKZBMrGlDlkAwVslkqMrGjO6xkU3e3aZyabRemB9fLwW5WJTpgmcSQ7e12Lt4Z
whjo7okKm49y8bMD0hh3lXPtleqi1MwK9a2ekltmoaK2k2eCuRa/EU0KijX8Ld9u
5mZzSqnFKofNEpS2SZrKaapyuauwf2dRnuZQsmLTX3p9YYdfLorqgaaD/bcx0YNK
REQ5cCyHavUABUO1AJJwJ6Yze6ws/amPKA4+vO/X6sKedMj6QTmMHPLhKzpViuip
3o1JQSSzKEdjknRPglruFQnqCRkgw8mBZeHYUuUW1m90hE1SjHh8Munsp76owDba
rhIGh9f1iuvOddsY70DhcZFb31aPavJj6vUMUsbulB3Za1LwYom8bGDl2POgE+SJ
T6CmZagKI+fJ26mAR2KZwteQDJgFxFZb6OBqaJJccstGMDXv8BXNxJ+wn0acHib0
pXkFN9eVnbp1WRDWSydAHUvGd53a+2u33fP2NiLFEhun1e/RHvCHAD/vANS1Xm0l
zHDvBJW/XF7VrutpMmia6QpnTpOs4uQOlj52ogMQbD2z0RBCpeqK8uy9gVihDm8b
lDXL8Xyb3IPYtkHA3/YQfAavt74oy9HGRr2+QOkRIkIcwPg9q+oOBkpGquBv7j5x
pEIdj3Z37imX/IzVbpMkb4vPaYIeSief0M8oWCxQOpHCeec4otqnEyizvWE5oK9s
TUt9LqoPvKdHXHelf0npgzfLWKnnxJfZ6Agf/fjeYs/bOjc+tWpTWXD147JS8pId
OmZjvsuKlJcfvR2bE7ZFgFhkhfprIxfBMvLOoxyLbk4i7RUauW+/KNKAcw2J0Z6J
NlNHG4xggwOJOUFVUB6JY+GF0NzjY8/ync2Z5OD5eAZUBFnsJocgazgobmnJt7ej
kiQPr2Dg7Ek10M1M6bxMw1Lpk9fCRspXvVzYCHg6tGNqiJWJ1GXabEDX2K8ilJcX
L+qZTgG2bCKLASbZHsUueJkJ+ZmTdm/Nd9PTGXKtJYeMOVQDW6R9e010F8oQsEMB
H9TgcSJyFRYNcRhu+F5shLsIBC0E/zl/bKCOdiYsrg/REIhbNza5qdtlpJPKq0J+
jq21SVV7F8Bb0k2SwzjOB5Nv1dBKlhgPeQOKq4giUuNoROjdSpq/YDxgTX1bKVB6
PlD0mDuq5IMq+DLyzjPI2krq15HYrntZCAR6Oy3enQDLFTO0Rmd3R8vZwAnmLqOW
D42t9upDQ/y+P6+GFZKIRUB+GVNWfjKOSU2dWWR4+V2CAs3vvCh1BacfQxwAYl9p
HjvPHYYFj/dHUQkA5ssjxDdwACvYZBeZMfjBl/cnzOZAXrhomRXYrVJsZzjIjBj8
l3jis4AR5cQy3K0Mkb+u9ccE8Giz+Vb0FCua9Ihx+a0xvgsprYnH4nnItcz29d4v
wFIt2OW5NBIpk6vNJi6GBBtG89xB0DGM2C7N6uHQiWgAiUccfkLqv5EECeQf9Q0g
f0pFTfUcqebzenQKDqJAV/oAaa6YwmOeORdjur9x2ehat3z1XFU6iU2XOk+UdVR8
dP4oXeYP1TFtQ1ZgON8J3FDeeYw/SnqhNtMvphccFyml2T9IpfCDMJWIrNxwPJ/m
k6ecMWU4Y+GSExDw07PU15/xUqjqCu1A6D2g0f+JKlvn6HoY4HP2Xls7H4LnovRx
5fQJ/cXrGiCDKRU+lyuERJRuZUT703XujxgujkENKSf54OXDncAbAsU7d8rO8mJa
DEG2015ZJUfDbGf1ZkiWnkOdpOdLYua3LIdHH6p0xERRb0U/GMRQ7c4gtmWeBpwV
aLq7go5phT3lIsQd3GBE13G9HWmqsF+8CrB4epbwht9O4yygsmSN5ddBvr+jg2cV
F5Zn5aDuu2yyHQTG2C0bz5mR8MwgCjl5eP8eqfcLiTCBsGiHP5ySAZwMapDptGo5
gFJy2MzeSvNvLOUZxo6eh1fYJ6/1kce8FNQ5N/VrUYaR9lPrnFWPv+Kut2VKF2zo
/LEe+doBJ5xgop/hHoY5KErTELevyakWM3IBovF42HpfvzbtItKm1SHUeQOxdKNo
OVGGUdwt7oj0eWcWdu1VIsHCDkP8j2DvpZlpdC31BsU1cGecqZejLGIfUQQYzraf
Er31iYWnsKIZbgQYiKn1p+uq677vYQ566Q6nCJRX9fs9xI/MO3/LBMC4j8LUVU3X
+kPp2pxhdBW6vLffnBFe0jCpSdhWEOnRIMQKfKRzWWtCEDAS86fkmyMroTsksF33
GnUoaEx+BQkDQlQeXqBrwobxlsP1cXKg5bZiEPScZTJCRH36ZWJJQnHgQwDBqTr4
rrQF4zHEpRVB+SgWL8nAvgAGRNJ6JXfsl8ANJdRv33b0wTNcwwA8KssLn/Y61+uk
5wfPySvFXspH+ZQm30a0zlRnw+7rTIIE9iAZzbkKjPYNB4NGYw/LZBK2JdEpGgNz
6Go8hWlehHxAKP50klGC8TTt5uREVMv0AZluWWQ228VL6HKzOd1pPoVinys7JkR+
7oyHNRpTwBzjz7v5DOHHuODlHDOFZ+9cskczPZoGxwIx5Oj0grg+UdMy7wiTOR+M
5Qgkr14OpT2DLiPN06Ux+lYkB+FfLMdGgOaMvZe7g03XWJT+8Nt4GZ5JvSuvUhje
ugETaJVRLAeN6UpMNuTp+RBKsEF16hkLJuHt8wbFDWdyFO3OGx/Yo4raSUdowqe6
Rp581IKDM0Z0ySfecUrJ9J+eGBgC2uwk5cGedYbX1SSgHkbglzgpRQeg++FmJaZb
sU6vhq/1gbu+lHERg8NOiSqKpN2C4nkk5t8+WVDG3okWmrk30e6WeeWe1cq8jsId
/wUO0kOB8uJglgl056J+4x7OYcM64Ils1ya1Yxt8CUxdcCP2hvdf0NG3Fck8YlBx
Lt8Lw4a+FuTWY0gsYXev5HzTOJho88OLcF5gyF/Cj2HbNh0pCd7HTNq+iqURVdZF
0cU7mCjWYFuvD3TEDw3E4TH4kXOCO0egWXlQeTMWUlIMrGyJ3BeK3TGDAQ/QjV5P
O8pwDz7biQmUw9XfWgqpV2Y1t0qKI56FQT0qjpWMunjEK7mNHyFyQ44vy2Wo1/q2
gDyXWqJQk+le9k9p9FP0KWV5xqAzrmZT+6QiAYK0he9YKHChSQW2D0DNWP0IPGhS
Opr115U1IsB9vK9Y8aQYUw2OvZ+AmsRichMGatZPcUG8dbRBFoxGAmK25HbOEjLM
MVCS+ZIhdMa0KKyVDl7b1BtGPlf6+VBfH0iw3VksYJsSCL8iRDV3a1j/0xjhhtSx
tEAmk4kHm0EPBcmciyv2pl4STohUWiT7Evl070thDkUwdAQzM2nDpsVEzJ37B6xY
LDE6ykiBIrPGliufFtduMkuUBIyI9uasTUqv8DlBrJZCz69tCtWJABzkRSz6RGe6
W+6VLTkKNIFGBDe+2AsCkwIqok69XI7PO7VtiLFLOehknCD10DKc3OxfChCe83Yu
iGJKuOEv7XMzBo6/gMQZq0b42K7qim7mHUMSQrlIAv+hQp2jIwLoj5vDQngg9lZq
sPbIrzA7oq4Ca/5XH7ortlkl/NS7XT+Vqr/gnrh4QvGDQe28f5mtZbBM1Mrxoxck
ztGFv88xIjKDq3CkySToWe1308DUrjD6AZjkD2sqwNTbivZQPKJk6j7dSMDoS3bp
IzQqn79LhuE6UDtQRWjiYj4CDwG/e1cN2YQ9fA3YXHBpq4HnNAZfgDTeshc/c/ym
7OKApjk959LbQ6Lqe5RVJaF69exuAIPEKShrVctkj3oZXPLZhjRapn+Y+jZQa+11
iymrGxSTRobKKo4cMIcMYKKVmiy2Fl8Rpk8SF38uLo5RSn0NICOYYA4HQC1J+D8E
lRfpDgd8i4dugs7A3fXvTVIdBq+N7pi6XDLSGHf4IKK8pLUMweZuyujsd0fsOlhi
LdBgVt4DCAQwpej9XqSXPZaRHipGbsd4LN4nO0LLptD8YwTPN0L2R3BVkGSPdWop
JjNKR68pUcc1RCAWlos7OU/83vqfJaaynLhonpgiqm8n1SIM4y5ivOrGMHpSa5/R
9dX1KSI/iBbZCxiapKBDxloza5Zw/Rb1N9SzmYD2Eeofw0nO710xurDpkeDp/VH4
g6WSysiv4LVqmc0QaueQRLRzrz/pBXMz7Q3PPIXbLpbHrH3554QQLAf/37GXFCLp
PxwlC4wXTO9qz6ZosiI04of4W+gX4lvD75FMqooD+gDEftOJpf/ynzq7FY9jO+To
eJHiJHprU9GakWGHSKsoHNGk1WMEud8QXRgTvfXLtrIZ9mAX2I1NTGXW9I4ipwdW
X0mT1Rszoac4tgcrYwouk38CP+3l6JhEuhfSE3aF1lD3Hivt1as+RO6jGlJZA+wK
Aj6y962tLN5sycLW8xBhaxDZbtUZqVNK7gvqpqpI2gXyVZYXAa18LaiQV4/U+bqK
SX/gNgru2TCeiRf+MVReEpo/qIkRI5cdEszSJ8lesQactpIGyhs8VEPHQXEYgXPS
NnL3EDhip/5N/DgBLguA3iDJIUePqruVlFkfORl/moY8/zH5p5T1ZqR6FevL/jIJ
Fgk6pAH35vvySwpqUn4RcuelFDwkbAHA75Rw1J0Hry7nkCNGMtvHUtNOgzhxmkQ4
ee/wPIuA1TfR7rIFVBwFkQikMvwJQmxoVpHtL31l/eam4k3F1+KdCoBZn6uvaNsd
8Uy2dgJTakIbSWNk+gsD04fsSN+LQOmH2XIEhsN7i7SeweMRX8eSMfPmZlAYrGdB
O0F/SQ+/7ZZAfbyOK4Fcfshuf0CVodfmIulzfljazmqOKWbsf8yxMvJ2/VgPR8uh
b/OV0TexQcn3y0BmNS7CvNKpXUP88eYsbZ1vkt0YNVJuhlaJZI2TwRmXkyP4WXIh
Iffqku2lS9sAP8gyg1sqJf7OA1HOujeFF/RYERRHPUeE4UUeJVkmAhbthqR0RPzi
5eh5BkyA4wmx4W9f0CbNREqePJCcb7BOkdVxM4Hb0aqpBk5bGPqOd2MfUGdPppH3
0vIOywLTFn82Vlv+n+0KRBkF9ocl9WfH2QPHRqvLYkCSE2Rtxc2RWmK/FVnGZ1ZD
vjEOXW5IhKevBJnWCKdYGDa7c41gFDPiZqT8N1Y734olbaRLFHUpO2midP2lZE0k
Khwh7qRPyZ+JXZ7wawylYqi6xxHJ1Zjb1WTFZy3KqFqJe6S18le9UVFTcoDXHNpx
y6hLnfW7uhIssDqTab7jPchKuZIJSzppMHZxJp8222O3FkUxkDdtlKMUpl5ZVfrZ
S+3bux5oCbPfk4jg5SCl3uZOImjnM4iytSWFU3rrP5fbEMK0121UJPP7doxFHSDu
yC0wf/t5xXYbt7zUvVM/U2m4RML2KTzsRj6mjOb4Vi/NUpBrxSuuiRWXOxWK74cH
Sb0ftuSUjSRujPV7iJyar1H0fhueaYuj1mfacbs1xqMjQpq3CySw2jK771horiLe
eD3aOKDogKSKXodhnYTVYVFAJLfKPdIcRTp/zjxOJZDK2bYWqUrBtKxGPcYkD9pj
SHpaFhFzJQOU/0GTJP5piEFM/AX/ItR6zwf9g+G9erU8tv974RlTbUKVq+la7uKF
UVKhWXkFtNJQfahRxFUfTCKrXv4yHgiI3ni8fJljRBRgmrpWEb3d3YP+bsm7yhI0
HL/GZdzMbEc/PWsaX8fFFzzdnGxhOUsiEMFhrV4Z9up8tBq8lgokGc+MimFzsLI6
4GobiC/yonAGYmQbwkZEEAbfmASGgpQy3OR45562wzBknIumyUKKz5BXjdzXVkM0
HdTlgNGgKUab8y/Ds0LEPTS/blIuHIKDWC7Om1zhozOZDSOrNXnyyDfvE/N+vYx8
vKfZuCDS4aKnFQ7ixwuA+vs7/usEAsn0f53m1reT5KcOR7PJrlGUvz3MLzzFJZV7
pAgc9Wz6jdQHfbv/tCCT10vNWV7OODIHpKhKtjd1Wu+3n+wQo6fss4f58DtGTn4l
Oi6kCisVjdyTaEV1AJTV83vAjlwZzHUTCXE2fq1KDI7Gl5dR3kvJuSws/5g9vOFx
9S8YwvXai9zIdL8HZnNt78oO2tjxy9Mupr7rZes5tGZvu1M0XN/BP7/O9tJ1n2A+
eDb+IUsCUqkqlO1+za88wMmQjLPaj+xGuSZv9HwFQPLOnPZaqKvy/Fe+kRk/4AWs
6bSbnK5VKVaOSP6lwyRo5Q67EMk0sWuRkp/I3FDR5XxSOsOBFXJ7K50IyJvxmIAV
C7i38m2jQ/K6BS9eLLn5HHOu/vUA7rJwUspK2hMCcg6emOCCw3p1cs4ecpZNk1P6
H1vGlHjmdn41wt/BU+EhsJ2qSsCqWXCcE/EYMw6vMv38q4r6lBaEMHs/fMJXD/6S
bxhLyF3seqW5CD2Vn6RBcxKGk6XCpdK9cTVa2PFwxUKNXH98u83CxU/7/AwQmbsd
EUKCR8b1gwjF5WZpt/Q7JooJ8uHkZY6NWXowu7e4m+VPnnSRdsqna3K+0RCWxUVJ
FRPN6/S8gP/c2P3sbGoo0twaBGhrDrLodvfQyud7wJI/L0fGd0MWAYug+9vQFjt7
jKxYicvGLQMcJHefCJnrCyhJdRCcJLy4kCoHJMKgXoBPYZgQdC4YNOx6oqR+AmH2
1CmkzAXYDTuuW5tqgIIp6kRxIDegM/qXic6TRfxZWwmzWG9tYSZratRzxDTTzTdF
oWosQKUskz2ANBlG1pe4FeUsqSjawFr/z3+ghGr5xYpXJOxm02YZXj9WHTCzUBQx
rCBjrIeQ2YUvKTvxN5FIz9ZAJRU1YiIl3xjQNSh6gy4i+GAxVHad11+wim/AUS6p
SfwYHANKI+Q8QrN0VTeyM9zPqwhAaabZZwu7mf9mzMoET/4SGggxfLXNVihbd8tf
ItTBZqcLeJYma5+4/G0Kw641Nhw0IbRyBkETQ2vxrHRuJspUtTgxkMY+clQ3Wxre
BIKGA6VDWBUiy0EepN7fD7fnYOJjMTYKCYUWubOxDkm0XEY743duLhtjO1HHlaRg
iqK85NfTsUAoOt+HBcdsC1JIyhWC1oFsDdQge1UcpLLYh1A7qqk5lOTWnPOz21sT
dGHHY7efqeV5dCNzituz25eWr0YU+7KFoRpufnSceZqIqSFUgT1G4Gs2VsTABkJd
dN/VgFVstnOl1zDMydcblIjuHF+tI5l7IUiF4N8Z/HI6oUrDeqg6E86kWxtQCYnV
h9QIKxf3VYZCOqdEXQylPN/g//BBky9kwT9uh1k5iPLsVGeyQQ0/ws44C7+1wfBX
RlRH5zyHfIE58KvdUL1ww9o3LYmb9ZDK6DgsGfA0w3RLETu003ijoDNgWGusUK0D
5iM1Rz/dPPsekEj9BN93/6+EBxAa3O8TIPwuspkkKmDvSwrZiJncqxhpVdNuAksB
Ij6Bg64YRhnU9IJihNhyCQojFL0tTXCqB51cHlbAA4KxeDmPs0qyz2AqeAUj7wKc
+U14WEM+pRaFrk4o+4SZwrOFQa1dyxkxRvx0/HWvGVL4yCXhfH+JxiRq8TpokDIq
IXnBro/Fbgr0dOTYE9J4bVhIphhYdq23Z/2eAJTHUX5umcjv9voWWttbcoFDFM3/
JfB4sMUohuATLneYzg8lIEIq3TIGcV7h9zMND6ps1aCvjv1g94N/jU/VCmWzlY6h
ok7oetp9VXNWge0eK1x8elgsHzqk2jOCjrbcYQxnP3bsUvac9nEc9+enyNn7tXZN
twLNnjO7U8vUGA+5nt51H3tdTpZD1DGVMDCPJIG6+8PNERr6AXvzrhB4larOXNTV
rpzkQ7RdHsK4weeO5AQzqD9/wH7tB7z0vzQ2Jm57isGRXFVpfzJ/WzF0nlzfc0dS
C+5hTxIiknXV3FFsAAd2SgBetUkLE0OeGN+CEYyeumiitvUl4Bhgc2qjBepwZxNx
ywpbn7xdBCZtvXaNnT9HwGpdrfH2Q5d48n888dz6LRqFthdFCup4Gh8pVbomGOng
15tGU1svUo5eC6ICbFGucg+BPBKHZjv//nyq4s+lBO61p174bSIhW61qvJFOCkDO
LCduZUFz6BOIx7gaOMrafBF3uiSUK2z+bGQ5Ncp98AgL/YMqx4R7Krnpl5GVftgs
sZNACVv5ORTA3bRpKHrt3bjz26DsrFK4H2IdCWyVBbdVuq3O8N/zG8/F30CUvKl3
ItGa6TFOwqSQbtfUcCICJDb0AvVvMrJCAxZ7W7ihjUqpqIIlLZgme0xlJBBN0oDt
w4ku0LkA5Ji1biUirumHud1fZ4k3hIs/yFDrfu+DhYcf96h6o+/7U0DPCPhwVwTa
WV9qGuTopPQaE7x7nHXUDLUYYOD0ryOoHY18l66OqkQKEUdz9MOCG0FNe6deNhbR
BzriIWM7NQzcktQfyLoUo/nfACj38aDzlDUXAKGRoOm580ZX2dpb2g5TM9F9HIUf
bFeBYmnE1+2P4xm29M1RPWcp3TVSLStdygc39qjWtF3DSMhmXyzkW71ESAysEa8P
nQ2DAy0y39B17+qeU7EYn5YLGf+zKbDiA3iX0WSYTYSfd6bJ7TfNxNeELYTCWP5D
n/ia2VaQFpXnr5vB984d7WRKD/AFAJfqZRIkV5t0i/xxPta3hZHff1yOnjUyq86u
GrKEYP1buAd3shn8rCrGM70CBKM7eQKKA/lYsCyR+o+Ymly9IAzLAwncCWXK0AnU
XQIOCGx3kr7esn5kAJQh3oDTkZ5xnQGZgjYyrHgYEaXSVlSEEOoqtvhVC5BdedaJ
Nwal9NZE9BGFojXLM2+g1i4rAYBhVuX5hRvRJ/Zs/aKWxv3VDPLKqGadu5KTf04a
OYEfBlBXnyUWZxl/UE7Mz2tklbbv7l+DBMNHBuzYVjah+rpUtLI88itB69fTeIh5
l+BRNd3K9zUe1d/9VMD9e8a5qux9864yYeBd5ww0J0Ob9CTSTJkjKuUwoia23eJK
h6hXNEh4rrlx84pdHaatJ7VDPvIqUwhkfIdUrTMuKVpJ687xoJrKbNoe4DAmnh1q
xHXEC4rBxdUOkc/3POIgr7O29h5dqfw2e3SepFgyHP82zLI6uqAOaf9VZ/rYciK7
+Znr/PIejaJbDwdmRHJycDfRNSpAvIJp+8/1p+az18I/4CiAt7ZMnUT1WiB42C74
8mfGUl2eFWvl+1I+EggiS/sm9j+zmXhn47jR27fQoSnz1BhmuOo81brcHX46j7lh
cngboGrh8ESFhLNkaQ07aAJ5FkMC/VaycYUrOsZHfRxt+G5g/a1ujVJDVbGMY/zA
jG5AO/MGT5quw8BPWNq/MNBwCgh1Y5Dvu0LdGFvGYwv/yJHBi+PpApYeCfx5RUup
GI3R6DKxpng05cA/rn0MxSZxXTLsqaOIbjcxYndZn7F1qniC6Rsr9J/44nLsRKIr
eVnogsvoiZROV6Bf03/sy5MV3Ch/yZcbfst1keFi4s3Jo1fHy7Mgw2cHvzMn7nb4
LkKLKSiFaCLd8EWuxZkBZKk9g48XIADzcko+HmhYMP7clPO2m7cwIwb9GgGVB66O
z8OZf8+HV6ru9VF3iwdRl/KAYb+xlzKRP3MHfl+C740XBjfiKzCS5ZnOMoxNNAtG
BdTHYoxYEFO8YEUB/PzLsz7z4WBu6guwsNzf7avIYSg01EfKu2gzXvT7JPsbjepI
zPxxuax5oMmgFO3CqDMFJ43qrhN3lYBDQfzVYGBE1NBKSIwC8ZeCD9kkTsOBs6ts
QAVMUcg7egYi1mtHpP6y31EKXnBYxjzOKM59LePVOjqLs02h/yAEv9rxtqbLRzI1
ll8GW3fFoCZ9o81OoXsKGHUvGaWas3u0M7eyAWhouIQLZ2rRSoGMg3iQ24efLmTC
0HhZzu9fWRCZtuH4e50U6HsxOg70btAeR40xcbSjRifr81td/qPmZ9GJh02msgTs
uO751ROP/5VpVV1MeVBP2i4JE6K9hZaReHdVGdd+ntylPTp7jqfU+x9U49pTDh1a
Iv9njKptzbz/SujgLJjqUH7+qsvMTc4sXSfdWDy/ozhBw34MkkrqnjI93o+K4MEI
07U2tfsR3Z72yA0PwchXzJzU8edE3WJd9I6QVmA2sPFSnQIsMUDeWgcEzYAzxNcY
USutl/cTfGSuJxDyJoOaTOGN6QDwhFovAOZhfxiRiVum6N94SQ2hoMPFrqexZbLZ
+Uh2qygj+jZaTuzxAWYtEXAQpLzDnO+9BXMG/JxdK8gSFtcOFo8FqxFpQeokucLe
B+r0/u+83mwYQvjvnxfYN+Rn7W8P7IS0uKdx1U0qd93Spv4RqDQZozwiAKsX2k8t
rmhe0s+AQBPpTkO+e48iaK3P6WUq6cloOyzdzRy2hNd9jGENUw4dFnw7HuNYWxPD
qhKviikSz/MN4jBhiicHmFBBZIug0JKLnRQKhxc7vNDeHdbE86C1W76/V8g0dXaG
SNKjhp4QixyrPP9+IDxXsQrOnyukZ/9DgSJTB5v5lyIdZeK/O9mpTZo5hTCnq1yJ
g/9AaHqSh+/7+5rmoIdEaBFtTbFcfwPi9d4FYdYlMvWxdnF+XcZ4xqhTrCttmaY8
UYtjukwIk84uHoGBi14+jD6ALMNLbLoy+vFJvCcfzdHG9QF/OXgcLi7efW4He+kR
32nljG4JrqeX6nQ7jp4tHeQ9fZEzlYRyUBKIbUvcg05FAHGRRY467JHAmxlku3l7
kGGDuhorhWctb3AMS9ToTSpGJyxLo9DqY4boBf0IolXiOk4ic5p5b0eJmv6gGJUu
VAwCweJPyXsyxMgb5OzxSDrgdyk5qB9318jwvKIveSnJsgHKZyB2F8pDQUb4hVCq
ZxilE0jRH7Hfkf8LmPx7HkYvAfKdaFwxVN/fUdXX3GJqItiR6Hs8WiWOprzKp/Fr
lJDF66P1dOXCiHhlGdYlN1SQatgxSjSPDcgcFwHUorPrJJ5LCCWd04B+E7p4pALs
+kBusbp9Mwvop2DBcgFtdllZxTmbnEvMabVs341xmiWN0cstlkjVSzrvyNRBSHGi
qx7ZJ54Oxz3dXHVKyDzHFkAdUKFejToXbAbX+V+OWLGNFGn09i1smQcOmIqUqXOb
jGISAB++URkpWK8Cpzj5QowW+P73x9mBAIMHz0HpL2Zb0+CQBWSGOh5DgBpYv1hG
gk2Ad4URmGcMTCtJHTI1ACQE3GkObbN7xwgTlRRAL7bpXQ09MJ5ooxT6wEpObR28
EVu7U9iUlFhRRmXy9kKahKa0ONYanofj2XaOWM9avsZXxH1hsrlmhn9u1l6VUcXW
rDBeJV76V7nYCdUEcZcgWaOWmTAfKUqkxCaTgPCFSNayK1DtdvfapUZDGJQaOCzp
p6sgo38/o17VbsxDvx/qxGfrfwGRkiEvoqNGq5WP43PwPnbUR32jQD49eflVvo8h
D+AjdF2LcRQ4J6JSoiVSqfkzkVuLNHgphaANoE1NxWSo/k1Lmawy6s4qWKxzu8y0
hJRNIaj4BcJvH5wkOg3DOPQPWDCIUP1HlhIIFuA8E67SMGy3bR64lPqR8C2Uwgre
0vx7M9a7UdBS1toiN15iDiKvEWvx6jwTND/zUX/ti2ShUxN0k+eYw6MBiz5KePwE
6B0PZguoszTwcxbDhE/WyxN18znNYivSJIKUlfbXutuD/4y5XDZ3z45fwJQC1a+x
7OsOwRtZUrWHT3NhuV02WmjLF99pYc/aPp4j0G7la3aJ/hkeYOFAfiD94aywrcvq
Z/VY2AFCFEZj4oDBiH660Ofd6uaLHfm4rdTY3EU5/LS40z0iEQCK9SBl+e7P6unm
e+/eo/eKphLhAL0oMtniPoFIPkrdluPmU7lcJ2sG3T45130KFn8ZtcqSXxJjmFXX
TA1I6yCAUbXYlaCBfWa1m3miEAFb0NoXZlkHzOblxR0BZKOnTdRDZRGTmdDTM9+y
hZ0zLu8AMHwmz3IybEyb9OVpFYEMUjdgf0ysKSbJt1qIu5ceZnT5EbMjKkJsRUlJ
Iwml2FFa0uNdr8lyh9TWHC3smCkpLnk5ZMUkcdgl6r/RyW/sRKUV1lZWD8RIstWd
MHAQ7ZlQMOH2z6hUFY4TpBUE1Z48wFMeuPbNpnwinMlavLGviqrbrJnpfrWg3C3l
bky0bqtnKLNGh4v3Owcoi25xLAeVIviYS6mUwCw/ZTYmgYwTqgj94nkKXcvth/vA
Pz+crEPGO01JW9kfwXVqkRAg/AGRUwdgP6WrDpScKO5lJwcJ2qMxbXLjSHI0YGf9
9YkkkdX/bYVjXgkF9jvSn1VF326pC2q1Uiy3eQQn5WMRZBHqE9Fbs/UDMO89cSCI
2FLymYQQtg7Ydt8+0qNESokK6VGfetTwz91ObNR0Y8TKHgsVjZQHlkstvXaUskpE
9VtC4azW4go5FM3AkuDUu0istgHi81KCycmwgVQg7x/zPrxAMLiODB2ajNinwKt5
Z8r/aZu+zsw/e32AZKaA6jOOUXT/wnKAn83EB27YjTjDq6WCJyRIC6tIGQ6bvPqB
T0CI5xckXWZmOTnMF71F2Y4eOgG0lo/B98BxUmAOzFGAt53I3efsQ0AyHY/eizGq
+XLA7NczUQVACQLaH6mkPHEUZjzrF1+PWGAwdMas+V9oEP1i02r4yxMCrNqvEagR
JzbdLcPBVxCiR26gWWhEThSEkyok+1oGoCNx2pseQ10gFKCnc4RcJ2hQVb22Felk
lSmhmFyj8WwNlozdDo8NWdhBG4j4u0UPykHe9jprjBGKuYmWX/R9uJ8IqGKmr4i1
pDOT7JyF0K8E+SUZ0UeOiSG9PyIQllK4RodSZ6zoSzA+2fqF/hH5rwm6mNwZKrx+
FC00Q8QFswf5Rko4YBKV/fvNBORUfJJOmU4mNaPN7YEZ7Z36udrShP0yzrPfFmDx
2ISVwdI2D9jGZd5ManNFGJWVc1Akthq3j/23BhQMkv1jDVlUmg/7NMmKBhNw5JP6
TugzpYfu1ANrFruZNOwsUN6kr++Z3mA8R/rrIJqLWdX1sgTNBtd80HjhnsO6lOsI
k7IXxRMDvsm8EFl8JNhm9FvAaykFBrjkuG9kXRQwDeD3x0i+3c+Q526CRJEnyg2J
FSYjVV1tf9ECTLgehM3rgOFUHdukZm6FoddgV6XFAOtT8j5OmOgp/ASYiC3CHL2n
+4BNMLoQsb3VIHcwTWDY/Q6dCbH27LL6nc7e+lr2BYxAnoabh+57YOegOIxnjkQ8
JuwMIARZDcaknpeLzLb5stXnRyT8lBEUmXWIofNRQ7VvY5B6set1ZQ/8WRcL4Bh9
cIwCcL2HxNF4KJ7RPDk5JSo7il6/eYOwc23fJa49GZz4sKOMXbVioXwEzn3uF7Bx
pVUV8hC1rVVEuTuNkMe+elh+GNohOI8MRN/6kUJfs2VmsNzJEQrwlOTkJNGq6Ies
7E1IV3c6xsRyFiBol5fvyz6gw9R53MZ+duMqww25TmAwusYheNGDC9GkY0+V3Qdh
iQaBGB7oDKlwCCDgXlPaUetqnnGaJ2fWWNXYHIXzytfdNedJpYfI96DpY9zKVMuX
m6jjeeSpNsMX0HOP8oNYz9zfUR04Ye9JKjAWEIqU8e/qF5wiEId54NTbor8D2fYO
q5+B2SIduOmUhDAAlrHb2jG4/OdC651pIjyZ043ZDKb3hy08Xqk+VSmhx2MnA3Ry
SoRsFdWi22BHI2UAJ0zdUA6rtBl8oqDcMdGQcedC6hStruD/KgaP1mwHpLOrwj6I
MrSWX7l8vy88s1ClKZ60QlSu69PZ1sIXz1AiIRtJDUUszWOBoYOQ4h5cHCube2gI
Wkfv45L2eFOk/aLGtW/nBaSO5drY9tKF+Wy8mYDB8iJ6LX/jhL6ZzF816rjJ4yN8
d7wcivJCyitxQOQPAxlg8g6vkUWqjrxBMzFC/vGUPXNg1yKcGYsmKZUdG7irGDyJ
jKVX4soYPh+mXHYK/ovGmD6lHTPZX3yo8ft6Jwtv8yJTPtOTOsfr1C/V6y7SwyLS
uZJGffAYLubSbuCaQskijJ1awk1tnWRCJmWKbPaQ3ngz22sKH9265TKcB2YF3dSN
PFCmxcEOGpFHg0J/NNdoNTLFHwo2l7u37uuCSOMZ+MrZH3E2qCeldjo54RunYO0K
5wBdnxFd5Rch2ty1H9frYFdyxAwadCcYWPbjnvta7wDmfjBDbaKWy5kmJuDuR+Bs
qo6JtP6wb7L+LGgyOpY4H2WJ+8MXLM5/YRwMYGTMyJA3lSm0fwd4TuzHf5S+XnYy
nfCZTTadNPvLG699Qgs5pdyG63UwSEJB2n6+e3N3Klr6hRufvz/1hcS+KY6qEw47
mp9yIRf5Z+RcTVdYgfL2SYjEB1EdaY9LvKhz0LacDZmSASSk0pidV+j8+B05OWPx
iivyobLzDO1MbSGpuGpYF5wiQJE/h6aqYE/ooEa78qrhQwuUR3DkV3SiRkLS2Fwl
i2eah5ss3BFuW7A1ebDbptYZvoH/z0uhqDf9YinrVuc/FTzpLJeg+1CQEZczxkfX
xN4yGx7Z3GHtM+/50F6bZ1FStds3f6o5YVMqqVi2ZobD5jDNvH7snOxgdADOAOFz
B8yZCHrE1g6Cy9LuNJcPCvfpmhram5V6I7zkr8BD5xmkFcWBiJddgSPhVSLLSOg0
VT2MZo0dGj+8dLnfHOYjVCKCq3vjnQ4eGGqr2E0Gv4WCA3iiGbCJf5EXVznnixIH
6/uubwsA4lOSJcPQ40l8kfB0KodrReM5Iuj5mPhtOFoZNQrJaScHpz8lOChUXa/y
E7rf6FPD5A55HVqstQVouYNOvfKbCS4YKvA1IjJ+LJ5oMypwdzUKAyvmxY9ygKXQ
s/wwddqCC/nr9jqZG73adt26tF8sJjRXMMWfjaiZRiks1BM3IPsFH48UnHsxaTLS
mpWNHu1x4YOjxQoalIGVi6Unhn0WbdiVjXmPVSqcUO+31roo1pLOyg/KoJ6Vtb94
UF7lI/JGtXtBrFY/0v2IscSWZpc2wGhY3a/9l74bBosaPmtSgdbwc54UvWLBFT3y
If1O4JvkvCFvCGZI7aaxhSwVOLOAs2is4YddWzCpR2ivkstCPeF0mE8Kd04CJRqT
B/areZTEPSIT+Cc1rZJvoqpSvbaAZBD8MRNHO0YUX8tyH+3wjm7bub8qbj79iy3l
s7MEOIbeNnc3vo3hFrdhtl+VA59H0tBKfPiL8vrPU2Yaj+17OS91vlGUP3b9QzAU
yHg4Owj+vDFLCLkDV/3Uk6f4OA119i/mNb6MkmBRnCmJiiFjSm3Cj5aBFwTTs/pX
jerq6WIHM7dRimuevqA1Fn3amK5SmuUB26XCWsy+oIkyaIp2IkyW8NRl79NIKu8H
9U3xy+T0DDNgaaLkcp3zE7m+YQMkhPdoFpIN2ILKCEb8Ttw+mwZraMLEc1dRX+vF
6/5grVmLQ399vUYMy+1Yaf08o6PYWiEMCpUcyBf8fdoBAbFlMgQduLPPh+17AIPs
ltpH3NZttPXrLO4megQu5CCTuxLJ493F+U9O4yZkDsiROanKJ0v++hpQdQzSPGl+
XZmTofJKIZ/Og7nhqay1RoPgOryCrMjTbE6zKN3yNj19voMa4E22O7+i10bX48Vt
piKTccgXbyXcXh5AVvGWQJrq+QEtCunRFYKoluMTmbmbRUD1MqmK7YwAL54cWih8
qUA9WsBoolGB5Uu61nGuU9vyWoLjzdPrvCiZNgJcxB0A5bBaBVBPW+wKb6IxTO/Y
WTMVEK+ewDh2iGX8BMNutIoBHEgb8/PxO+BAwfEGYepGIl+VdZxyjuE15NSzF7BH
czNM2800E/wvMZAk1yNWfk24WukadwFFub9BcDr6oNiQwliKIx7JpK7G/dE1HQaD
a4XxekWIodUejvzARrOk/GsuahvddT874oP7L6BEbH3VcUy0H95YlRiHp7ExnOgV
3H92qSFVBx/OHU7RmPFoIpJnJgbgEo8JgRP8OwbKRC7TOFs8DnVouSv0FW5qYI80
s4j/2NoFDM274kJTPd/mixFYNVk/5HZh9TJ6OIGi6z40SHpkpK5Ck66yWzoSGK+e
/vOQoDiQ2ItJu1QsevF+avshb+1SQCYtRXdkk3M21Uo7mxG6ay1F/EcX/7GKZdms
sWXqb3utC5+ttoGfU2p0Y9LGfyn1frb9V8qyjG0GGz0u4Ml0kGU6yaI29ypXSKLh
QqbhrMXnFWrkOpn1GBI5Ef5JcR5O/y0wvmBNyVV3bUSQCj9I7yHA6oYWR58WTZk+
ztMxOMbnUHQtNrS2N4Amib99dAM1Ivnqz0NItwUUM89/PWoBeiUpfX2SuU80JYmy
OCXLGI77ZCRsOgUdEzlNtaxohaQKmj3eR5xYdSP/UqwstsqweuMzIrAZg8xE1uyb
70I/Zkisuf2dkmhAx4mZPA7Pmy0EaZz5s/TxxJsUdwYxVKOtUPtvcUdSIqkMA2j3
p2IFTugYEdaiZeGpbjejF3qQ1AfHLi2v4q2ToTHVbe+oZL4+HSF8g97MvJhLpfDm
uTNWJ87DqmzzYk/C6tLUhctB8opDqrAGmfG4RWConwSi7ODivS0x53kXckWj4j9e
G4DSOZzEK+ObXNCm6tw7xzSm11AFumER7EJhB4mCnta1mVerO0+0Pz8Z6DxmMNxy
lgSCg2Z2Q2/SDhToOvpHXj7WDTpwixd9KxvGwz1zoR6bbewasvjR5x1QXNh63oTN
uqb5Z5t4pe2pl3dOh7ACEkQW3tKLrgNYeZYuXqeGMRVJQYPi04+mjpkNoyUsyP/x
E0vUEn8qoTDK/UskNAvcq6J2raCaxkkkUBkNlHOmUzGL80Bc54Bl7AxBpJg7fRdm
mKLJYrBks0jEcjoy+f7ktpCyMZjO9w04vG6fMqjvxDRpQgI1bv5SOf7LvFlSu1vz
jR6iGs3EHeGkzn2erkVi7Bi4azssZmlxwWRHjVIIV+H3W9CVMXyrMb2jEgiTNvMH
bi07FQCuQMR9H6n2eWNXaBD1q+2+QinyU5kPDcdv9phPJ+df690mxrKnud3y+tyF
UTYIu9mQINbhfeLBnhfjhzmnlSHi+CzUFcx9o+ByuNYE60X5oghKZopoSCDjmcim
0MMWBXvX2zay+ql6MqWbuCLve/O0EJ21fH+p8dL8uDNHjR7YV1nMMS8TWBUGbKtP
bCpmOBEvilNXis/YGHRJBbzAlqZAxwc+RJU94PvGAhIe7g2+4ljvr5pTzf28XKKY
fRri3XGS5ZV8Cu69wE/qiU3OmIzyBuJ5Ew9aA8UslDLT8rq7xqVgwwtKT6jVMBmp
HeQeg1LXYsJkhKPkyxnt9xp5M+VloEfuYd7tfAOP0D036K4OjzlPHGuhrMSNfB1O
ak+jT1KSJyoiGEGyulBQoig6NCbmTNGsW8PfapL3k2RlZT5Gw0CESsslX/aV0EWM
z5278TdY05TYvVSb8D7vzL5acEE87nOcNduTUd+TMprRuMRPYRPbNaplq/c3RGWi
Sd6tIB+yT8UXevh/JYSDVrJsMSjVHiFVliI+k1Nf6Fc6aRwCkLv17BafMsRB/jt/
Vz1V13RIF8eeTU7k+IGCqCoBV3W4UqIE1EsLdH/rystOmabJSidgco1dFeueZjlD
ysZfJv2DxxGrg7Bo5mgMUakp4ay5hmD2Um5kRukIkIqEBePJW/b/U/yq3Ufl46xs
Czlx9s7/+BUmClHwI9A/09w5OUsl8HUNwRuL87KmTJ4EDqEFtOVZ7AUAoxZns/la
CPdzTQzNrkS1eQnz0WmSNKhKlekhRQ0afB36th12o6WmzhHLkyHfEqGPwgLW4odG
WNPHZdKcSYi02ZIVDK+MBF01siQfjF2iKNAmtKyK9ByguUUTV9lFghPZg5nRQY+D
wJlNyex6FJt95UXwoEldAtGSdntXmgZpgtMcZWxACtEjH1f/Qw+WtqIkOZS7uaUR
josZuUa7eYmSk4/55bkBXLO8GNNYwaSHebCP8MAejSjQH1EQb/6BJI7WIWCTEyPQ
d9EOZJE9oCL69tANxrgpExqhX6to4hos/E1KZWHKGCvY/4FUAUWkgh1a13zH44dx
qrJoY3Ipgn45smmkZ8TTHszFxGd0CZOS4qi34CUXtxpQRgsLouCrHxBIeqndw1YK
dbz9eXgn5YCBrDwDXN1zJ0qlnlLpy9I8zm0CCr8n3hZjlm7H5aSmFgNTGxOBf4BG
Jm4XG2DrRYy02sUUK7OjPSoo97nyV8YPgTo1WQ7ujLnPQPu918kIhzN9jyZUIZ+y
QQAkyY//AS69JxgwVL84edFkP3KqMsfkfIRtPOLRZoX3gU4CXD43rkYAVUTBPQSE
5g4cYSskchAH9kXvCnkiru/FFEoTEbEJkf+2M107rS5xuzUMy9tH9rL6tNvsQZWv
tpRRYqUIAAv7Umukcq2FOqR1ewh07XLQHxHx/pzFz7S6qDvWo0JOe1xxDRpvr2qf
2NXoALUfRyKqcnUuYXo2KjPKVU92EVI0RsmnnD/SY63BIxqE1Dtmup7Xu+T0oABz
vAa1khovqA5yXuYoh3efkE40rQUABcFuoige48XkS9ntNAUCU8DTncLcDsrueTPK
CdeJFzcdtz2Bu96txXnOsn4RqGf456JP7tn3PbMw8Moy0BoHMhAX9OxUWeAEgS2w
XmvEb3TWHWh6S217H4+dJLbwncanGZlRCBdRhRoQbYIoIa5g/0ln5GXLpzciNwWC
IDCnIHbLOPtJ2aIxfgqXyK7y+dAUaDn2yjc43/oRvvd3ivOoQnkRL9WtFYtC23go
iv2TSnpcINE8Lg3MisvlaOJSN3nvO7SwXiJBZfJWHLpOAsVShwziDn77dLSeV/GX
XEsTOfiBjLG05X2Izf2c2ID55eFj6apx9FxNZEIm8XhxyLm2J/BzU3pPgoZdiUsI
+O9BYYoDoESN7aBH7aKLMazbWw8cvYRHidP+GS6J65o4uqyQ84HyoJUL2KT7Ghar
Nag27OnH3qSRy2VSn+hr1PVqAynmNnYNNTSZFMyMs3SSsPUA6GDHxLPX443dWPWx
KMEz1JvaRBencwpEaLrceDzUvdACPcDPnqLccZG5c5Jc+o/Wf5azcokrlkXpqRPh
bWFQppx/8dBlGfuybBVFIHh40r29bn+NBpkkO18irrIEOtKKuV4+cbq74pQnqI7S
MxfK+SdmN2vwQj/eyA27FNjiMmYYmWSnh+rKYyuKt+ETG/is18AWdlvxhfgTDjvY
cF4VdrR+WE/DuxssoJSS4K/RrbAZmoYZjHAefiQYejIUrW2UltmntvSLnD3P0YsH
P6o1sXmTTJxocYPXt6jfjfADeNwjYF6EQuPX5b1rAwhs0fNvT7im/KC85dfrUyn4
ilCzax1DsQrn1tWKrRQ3e20CDpmAfwTUIWMy/wVLf38joa7BNkiHpo5tm23Oo0Zi
ikktha31nwJHinmUPJhjCt/HlVp51z6oXefwy+XyXPuW3/wATewE+zggoKxyCxAG
R2WMaia5vEAFIxAqdEt9VIm8R6ECY9glZ5HFPDeeR9FDa05j4a1NEvQ+DdAQs5qB
UsTA7vwxmzvb6apMQ7g+lb/autO+ILGTkfGzhDc3tNVTgWGURbdUUCYI4BKYMwwn
LpvOIvrvsryER9T6nixry4EPF5WQM1mor7m0biHBFTxjEpDiWtiscf9mV3X2HV70
ZWnLcyWIoHFIOPql9cwY9KyTjpLwVQgaPdJJ3W8cas7QnZ6enKAyGUjuidiz0FkH
UY7ofWStVlb1jyX0QYMiUQCJSudzy4/IlYBoUgPl6404G04jDmv5fTL7uNxuEeiv
jZ2m7krnMhi8BZ1UFAA+mgpyv33qbD1hEFIc3Ph8kDY074n/18xaD+djXkZY8z+n
6WlA+7aikU2zt7SjKvJovjiFqKo/vfLpHTsUyIj/HmVTmiYk5gRZZ7uZg/7pu7EU
8YbzSYXwUia3HSa/nUhzOT3ucK6aBjtlEfU0AqfISxBZrHpDljmk+BNqaoCj2C7/
r2sXFj2iJYVyOxvfeFlwc35CxyWW7krU2fOuZE2Ro1D5ItC7q6R9opgk6blRdsAP
0HG7mDwUqyb5EAYgY5c3ebD+DAP1fLVJ/UEPrG81D0fCXKzD5LOgEGh6iiLc/a8q
nc+Covs5yZNeLaJIL/2aMJb/9ldTCkRa+xaXR45nNnGoQhMQAKM2u84QXRq9etxz
McAamsKC8lbFeDh6t1aEfNUp0vIlZuW03xVsttu0zVzxycNDet2Cb3Qedf4ffVcV
qqLb1CexgYRFub4lPBxtz4DO+ijtD45SvY7YfjvCnQibwCD6xeUTcEww88PVFla4
pcWtzrF0i2665WDKk0JWmyA98Tb+sppvVEfGj/d4bFY0mv13uo+3UlztP0pKCTAa
/hEcJolDGzoolJ4aKVNwyF1Px2ojHAiQI0ztT82KMrYthxzapfWv7S2Bg+D24fZU
GZc8OXUJXUC2MfVmrnSc9wSHE5fpypj+8/8yPfJj1L43wtbkMziTxGzJvIvih7IG
BFPSt/r4vb9VUI2Q39Ocn889h0UiB+KJyEjttXsSsXlZ5T10wqxlOD48a+xIKBHT
cx4ZI17UJ6kuLpeip6cOLQbmFECi4hyY+gnaGMUf4IsMxL236kCamvkpjv2vp2dm
B1CMZgelTEbUEI723AwOlMxmGLIGJHIFjQ5pCZ7rv3JJM8dafDpW/FRxNPEkKNAd
YUs37DuI8O1BmZ6xCuJ8KLhDsKXLTpepPvo5VmJY9L8cxBrQbOEIYVIoj0QEufTP
8qnJGGlqTgB17PRt2mMvytFil3Le/74GOmJXwP1ads6WL/I+lRKMn44WeoJeF4Qv
+fX9VcUWrMojmBp4boMjnQHHdZepMHTqYE83H/zxmo95ZhORa/MVRICBQAq+l5c+
JKaOEXWV+m+ktZuzn4aDgJI4lqqLuOm57kQpE/OkAy1MvT0t6kYzoDmXvh0cb7El
Hwrg2qpkc1OUyv9CoRBqkT7Na7DqPSVsXZCkTsCbZ/Zl4ZLDEHBuzHBQBYKZ8wiv
crPkr6DoWE7mqByKTfgDutNukNkNtzuacGhDZt2pztyyz11fsdcX7s8KZZ4MkKxY
qG68w9RTvTK24sg7maLmL2BJOAY0peAZlwRKKvzgVsRPbTR1IcF4glhEMV7eeiNS
VzjE7rAZCiJB2IKlNPKMEVUgoQxbP9sZJIQyNUZAVc9dUBxORxf0A1G2YDfm300G
279YfiOL/t1xaiWAAOdHSIl45aQNvuRGWvDcjLSUnYjxDWD71ZH+UDMYONcygTCL
9a3o1id6WDaKOcTymJp8xJbM1oN7f53Zbnmk69OAkk/V1BifIyLLxFtAIw5zMfmn
jw7UtF4qMnAMp9QqD1X4nhQS/KhDtFLNsu9k+WD9TSHEj9p2VH9B+QjQPQZV5Rs3
uPm8QSfibtpfphFV7CkNLeXT6+fpk9qdui5p6NHHf0xhfnDXLPxQDHZ7rfrcFW/e
YsiukBHn402iGQy2DPpbkZz/D3F76LmKjTJxkVshccvJOy9LyY06Fd4hJfMrcWey
rakIMpSuFRM2BdD0HWavy1hv1j1D2aIaZPcKKsAGB9JS+Tl1yzgXWIR4pz08D3Aa
zvfGj1OA23f23EbIdKCcAAW9f87QrFzU6d1EqwC79cKSDzAExp95w0EXxVJ00C2P
xZ8ok250tqaDpAueTCHgeu5BWykS7+iRnYUBkUCgv7OCwmB2aQadWOSIn4x93EY2
TdMUZ1QB9Tnp0p+EBAI2UqK36/Scd6S01aekMqIlywHoTRX5Y2107wzP2+gsKonh
dXvx8HsVKahXeh1Wb2GHmK1zEitTYBIcoJriQb22EdQ1+iPYsRTOzer43H6e8deQ
4e27vPb7P4YHh+lALZYrO07qupKyumRbVAQAoPB1oJ28/fGjZUUyESRJqeBo3eYb
t/78ElI/5+HAaYRA/ShliCpyQn4vpf65/+b6BqtSGAoHnA/So/4OoXwHlbLpsDYf
IaF4zJFOffjDMciTdsUgmgLkbVKtl7j9CxOl4SuQSb0+d7kj4Oa8/yXHo/YvDuj9
rxq+NYgXyzrJBSWWo0Y/K22wphneQ95vDy38IwvdDwNXaeS603Gh2l05FIEosdCz
6l58VEguzBBHcJwgRavZ9Waim3z/eK2QqxET+suThXJunxmqPm+osrpfVvry2gFQ
hHVK5WxkUigrAS0MisVSowB8iFA+ACXudNjkpSBLmFUCXQEfOrLurtRteDbPiFFp
nWeejQPt+9CJwgKOLjJspfC3sKRBD8DP81Hl5O8oK4mfU7i9PMy1lDrZrRxOvhdr
iFgDIbg+/aOG2L/Xaa4PNdrooowzxu2quNnNv3A4c+mM4atWaFYc1d+rqUdnnF4q
c/ED1mSe4HY983XtgbhRrds5YEysD2D5Ypn62ksTByWHmQrmVgXkhqFsDpXQE+jx
opetI4hW0Ete5qY9Kb8zXIWqZG2W3mMXcLC/w01M4QnYjWH9e5S9yb/RXBD+3e9j
tvtQrM72C1h+7OgOwUj2B/a7/xAx76iDuxt3mBAE52RuBVaPVXBskQfopNSUsrRG
Cussa/RAUvmxTIlVlTr1b9F0FhEqxYgt3TvAtPuFHPhn/uZn0bOmTC20slNNqR0Y
CKfJYWska2gPJQuqWEsI9uu6UuAWiN25hbgwho4Fsp00WyoOb7e6V2YTaIejV8US
VRTBuZh46sics7eZRvlAQuna8ySsX+As2ZU88nPCzdl2P7/+8Fczq8gxArhGWSEE
GoY7W+75Ff81TMatsST7Qau3iQ4ZEY+sWlPrtGoIlXqOYD7LY2Qfh8DYuYQ/YRTp
y4siJXasbtNG/J4G1gxDeejOc+Ypo+ERHyT+5Ybf5T1By0pTyLSMv7MAhgleQsaN
+LuDqVIbtYBW+8WE5pLRLTv0jHM5OcmXdUgoFzG6/m1dk5Fm6jogeKo1yLQrwe6y
V8J6JL/2A6OextTfOUZGXSz4TiXNe0cVdQE5h99QHoII6Gr88qEkBFIL416NCnGB
VUdc3yHBlGH+jjPGF/ls4ZsBGeoy9PpT1ft6TBkVMABUN5xluPvdEFlFJR2kSFK3
FvwQ/bhMLnqt1YXcl9YB1Jzbzju3bg/C3bYrWD8L1UEoWkn5Ns5RbOYqhVRg9/TM
cLl1y1/n2twMYs/fj9ij7yDZmixofiGyuDMfyRTowKDCYey/WWuxLTjXE7XeD4+I
Ii8X/fRMwG2+exdWoLVmVOzQFsn0hi+Z5irOmID3lfXhogQ+T50y7o5AcqTpzZNF
P0WQJPjjsnWToPesX7nikfEHx482vQep/koSBOsIaoH90LUL3wQGYTtbcynvkeS2
T58DTU5ejo0OS8Phc6YcLXtgFvC+ZfwKefuA8gMJc2ULkfKMvBdMj1mxDtPfguT3
notdyJJXk5MFXuNSe6g4Zaey+3JvsSUcvSyhXGp9bw1/+gKe/cDLTWpiCJodwt/S
j+Ss2X0o0QZ5Ix5xDvvligeowDy+7MSoBaKz3AP55F2dW9g5N+6yP2m1r6o+7sX6
XR6vFJi6PHhwKj5WNjowNN/ORyphRzdfpiieNYe1hEbu98s65uLPfRkV+3Ajenhj
5FXV2VC2WVEo9l1mYYRDqcjlIUVaTr6vIHT+cg0IP0Kz9GVV3WwRZwtA73Bwpnb1
6owZOMvTobpULH5oVw+YZ8e/7pJu1ONYQaVZM/cUGl7WEhwXm6LDrx3Gjpm3GPV7
aN7FIcN6cg0o6g9mU+gC6XpdRbejhWR+pTDrUFiwSJXC8PDY6bxB/Y4izvYnBPLZ
KYfYmNxb4vBKN1dWuFJNT7dlmlCm3kaI7IoM5Bbi71T1b9eScICj1Tc/Ec7JWW6o
IPfTjVRfjciT4YbDKHXRFgBfGcpfaQXrXNx/K9EJoajO/vfDs7fjLR4rZRf+0HrI
rv5+YYK8kXousnwMjS5ZE6SBVb13ztPTyd7zllQ9scmTxNHy2NsD3TXHojvpROEE
NhExdAlDvDOyOCvtBXmQXMI97x4zXCJvzOAF/QfUkoKMADCndWK7hd1WMODEHC6a
N7a7IGRNN1yiMJHyf7OG3n3FaMY1XdRPsuGlWztjaw+H21WWjmUBFgfVhMbeWqtI
AvA9Ya8tRQpcdirt/ELCOs1AnKodLJyuE7gYWm1mN4UD6n0myA3Xxft/JDvXo3lw
f84PLUMJtmIzTYy1cNnS6K7Gd8EePTlXfFJVk8wqpJRXLhjBKs9YTv8Aq9XbTcJd
blRNDKSwUutKLH0ap+Nm1uuscokm0C2WgB/JsLe0dFG9w9RipHr1DG+iAojvJt5G
Q3SBReP1n7XRboKGq2JeFP/0rdXh7BypexHDNy1vLIJ+5+2h1AEwbpkhPK4y++pW
CzM+Jwcbh0xcPjZulMLaxzX0NfryPKCQZX2dBv7xz3vxzycrZlutgxTis/bSiyAi
m6n4wdiwk41x7+5Eqy0Mj3xT+wZKUHid3DDXhce6R+YxkVa2k6qGGT17+v2g6oC9
Un0YTmaGF/taCPXpUZGB7cf052hnJhTW6CydkeCsHYz6QP9M2kqa2GDweHoGbEiT
laz47x1VIon1isYHNedCiAg/WgKP66kN69WU7lWjLRq74OmKwqfGy/bNjxgC0z8W
nGshJxu6KjB2aoL5+1x2n9PbfuemBeHoejq84RTC/OazDkaCjg4Iqs3/wawwUVvZ
YMyi1tD8gTzmshggcPs+SGRzQvcJYzbRpnKf5UZofe8FUvLLN8EW1z5cnaBjEbWu
/e8ll3QRqFiL6Iu8zTMDmrbWBHI42F2Pz44JBfyJp1UpnhECDP91m4c+t2l/wquq
zCZR+d4w1OJGtS8DNv08YfOzTtkrIfbt2b3+bnsOTkH1sLvI9ndv4AXcY3OAIx+0
VlxcqRod3s/MhZnnrUh+JGBpLY0QGuHjfNJgUzX3m5u7r7LYgeQa8Hy5XLr98UFK
NbklIkqozR20EkrR7VQhLuxrrGP31kiZgvCNPW1JKJzChgfNXnyvb2NlbVUUAMsR
SdNTyq7mxmZ8Vi485/7A0TJh251+EnM/Rwao2Kt2kRnD6Sr/ghH0dl8n6QyPJkLh
GZvifMVicttY5sAAsx2jfDVZYhj5c/znA1pjhwF0lHS5Dttw3zcQMvHLb3ad3D+j
88vSpHA9wt9Igpr9SJ/JZfuZtvcRWOiod4wDWlNvOTEaa4REB21yhXkRJjMEpnpV
2kn7Ow8csqGOPiEKoH695+99mfTffzoxe+N0zHenlFBdx4MXGkWt0Bvojff5bVPU
agBdM8fXQuMA2RKBKLX0tvo8CmhPZVvDHqwxf9AOx5q/jm9U3nJHcsjhevY60XSp
8P8Rmmc9SF7SDYvpocXgMc3pd0CGWyz1ExAmxJ0ohbkVdHXsdHZwoK5onDGXvkdk
zQVAKcf6Pt567Xm1vr7egGeUK7o/tuX4EyCyg6c4+GAof+x0WesTLPiedhZrfAaI
FjfQUzIsJyz10nwaAeFWK34Pz1jf0TZmVuZ28MlHE2rhhDC0xNU4rRMVubNId81v
Fp1H+9M9itOK+rRbZPokwvj+euRbI6RqXUtLOwerZI0ynEzo7HRJ3Hxfqs3s9Oft
udmEtBQr5geNE9cWJIvT4HmBx6R/BKRk7BOjcpsxeK3xhJDeZp3M82fPjiXEAPGy
qnWfHEVRCFk7buxHe8YiGY9DCdSvzXk/IcXjf6BW3e50uhnfvd9ueVUvzKeLtcZW
kWvTCCgD1ueBZj0FcXVpvIBqRZ4NbXknapkI1OT98xBOlddLzHV1wzhxVS5PJeB5
1Eo+s/U0Bc3Hllt71RuKrmmBuScQ7GUK+cQhwJCo/udXSK6LYbTrlrpPcvzaD3HH
wcmUviQTdhHiIw40lsGcHjbmn8ktcPYQdTJGXFW4pUQCZ8gZ+jkExHXKzo9UemHr
Upg3RZU+C5n2c9vKkX7CPY1ivfluKFBOMiDpaxutP7JgMrUEmNAb5JtNu9xoQD/o
o9tuoJom/ouLwbtm5poVaf+Y4bZy79WvkNB3TmVUWsUD+odo0UslkCbPTQ1yv4/l
BXn2uu33lMFUqcx4cEO9PAUR3oPG85eSovK0UAFHjaRCoHXHlo16MUQt8bJNTTm+
+iPpYmSEVHflpyJ3h+GT03A+tYL2aV5arEO5umeaAfQTjRxiahveS2RSUAiaD4SN
X7Zt1j8nOBTiPpPIf1vlxhPmgrbvPdsOtEXqXwz20TTDOz0I8Z3I2Ya6ZbHCvyxf
ToP7c1G8zjv2OgUi4Vl1oyyyd4Sx9Twpvp8LtuhecRKkJ9g1K9tYSP0jsoewpDJI
UQUUi+PwM+xS7h38RU8hAlLP/LehBOT4oAY4lx5aXXN6TVABalP8uvY/PApAuthn
26HBecEVoruwrIJhYMb1sLREjwT2bzvHDsOAtIYt+Huubyo0kkIlQGJN6D4IOwJj
lW/0q9CLm8Tsmea2jcHv93ZNkLcLC+24UGgZlqynAXiTF5k4qTtVxiu8J2Mdbgae
KFTNXppq+rR+NnNIS9JnIW94vVMCj/ZSXgyVi3qSgZnPHzqDyzCCnegpr/0boo3g
hWz3VSCMw6veRkiz4MLvJKKs9e2JuxWbcKSb5VDfcxG2ziunws/7KGsWbnzV1cuI
xy8wENwVX7l2x0woJ/MGi5C464Ky9jDyAnelASBJDo7WpdwlW+pXymvibMu6Zhws
wrgylRfaSK3hVpa20pdZxOh+JKSZDT3wcEOipdojYc1RROTwMn9383LXxuGU9AcQ
aKTd6SuIj3S7Ueb7iMhLNX2SEITc/U/wHD8YSkf/gpGl7zeJUQIHliPhkZIHbfe+
G4UJoBr+129Xpl+P2AeMftIdcwtoCBXJ/VWeOopKPYm3WgUWX0P7vFgJ92pEoFqD
rDk2M2K2Fped82EQrKvsMmxFGWrl/OAAqVTdwWre8M48XqEv292bVv33kOnaVle4
7QJx8NOwnfUraVPOkAHaQtetvQoLkksapkK/9HSjvOJCqIcxR2NsykaKOZvdZ+BQ
hfvBCuFWrMyUxDd4NBZo1guYjl5pa3AVRnWJbBOpr4i+luGLGf4+MYUoxoLN5MRw
MIx1bt0fdFz27T3UEbE3MXggvEl9+otczVEgPpAKRPggeo+FhIsIP3eOzCCf6BAT
N+qtzLNbPPjpY1OdsA1mQsQWhTN+OGuunvnmia75aCM/x1MzJqmP5jtj3ahquFiM
b4G/XxpdMzJ2VShqEXBCw0J63NYqQb2XfsyEfUArAJIfUjDS5y174qZxzgVWe5Aa
6LT+PP8JUbYfHsXDG0zD78TkTIQacd53iAltWlw70Lh0dNv4Cxm+fDck5370EPmy
A3WWI++DZmy++vHAzcIuAf+XoJZ7LzZAmbfEylREiuX7uAq/hSNaJHMP/loJNKyd
jZmZIa/k4Et9gsu/B/VAt0a5sVKhLEr5VerONjq937UcYxUTCXhl8w6PUwblCZO8
k03CcyIBmFilQ/2H2P3m5gShfC657f0+SUXYV2ROsx1DpdT17qdavo8Xtf69U/AN
vAk85OWturlt24YsA4jHHbPo892JOc1ucTYLRozMahej1JezKuaaiGJCJlOsgxe3
su10jVJXFCPZdATbX1iwSqQ/HW77LJfS6g+F7WvezbjGcl0NTdc/8YO9gn1Wxr7r
vFUqrXCCAxBNU/GHKUjhsDYIkERoKtRJorQjBmzVJ0g9OKzn4bUv8lwErabYFYxh
xeoKiPpvPQSGVOKkbb4ajbWCcs982BHQD5B14j9jzNSucMMG4088bYSfnyRvCeJn
Q8VvKa6juCxkx8jvgTTz1p5fQZkNC3L+GGNIH+1TlBj0zrR8naee9/T2yfPz3wt4
YtswMssQo7098+qbyWAz33RY/0njTypXLAPpInExS7ZXAq+u6fVeI4wYYTUeZJSu
u2cvu0zW4zpJT5Dhx6QL2e7YAh3jUKsD5mKEP2OC6iQjkbNddJ0p2xJVCBsqURC7
bpHDq9IYXrZPfq3JlqjxE7c/PO4iyViE6GMXL4lwrfFgrcACWDBxqqq7LeHdK8Bk
u4MkaNQDxHBLcf/vGtNUSN4oH09Ww8Hi8EV/ibjV/KT6t7X0KERVMs/0LpPLMpDq
TMTAIvpQje+2W4givzm/QtoCAY1potjQujq24xHUkic+Zxnxi01BZczXbGrC4+2j
CB09+/qFo1/LM60V7gwZfXQUc8jfAE1uufpcIytH2vTb0bmWKT96Cdch30R8PJtw
K73TqWjdiqEawr2AJf4Oy9UfyefBJ2PtdD08rvw1STpOcOeNmWKfrKmpAqZ6f7E/
qCLmHOm74UEsUyjd+lwGY4t3XK1rgfYLhgQi30MIG6cK+mAbmbKXvCKINSOkyfS+
UIJmWf3YwVKjIXy/2zOV7prPb+A9fMq8Q4/nDRcziZmuBxtfa2wkskuzaOYLxktw
Y4gA566ZUzxFI+je+DCAPI9vCFfl2sVd8HUgN/YKlbl0qVnfhTzivejzak3S1agJ
9pbXLhBIwdzX46xu2FRa10euIovJyIsURm8cn7pVHnjBOS4JvQLQczBhj8JTEcR1
cAtdoisyYFkbwS2jOy1bg8E3SYjArdLV5xaJow3uNrKkl5qdqUJXVatI1pTMD0Fg
8H89hA0cIi8ITWbZ3nU5IlXEYz0xKlwfA2rCijUAyAb9hwZ6y6sYVskmEwv1MptR
ZRvVmd0vY/5lnAkb+Hk8VmvkYLBr/YdR+69yT4vzyXFyh0DVSIMLhLbDFLYitl4v
TIXpP4cXvNo7u1lMzAm6mlCFR1Kq0doJ3sdCjJcQUGa/jifhNwh8w/vocqP9P//I
WaXsd9mPRGVEPPE1BVxo8rRMdte/p5+txSNk/Z4tof6u5FXhKg3lvqaY9wgsTwcT
OapfRYFGVQwHN4FU88xKAYkQ/NzRcd86hNMnOZwht+PYdqXsPIeEshtbVITsixjR
33a4e4p59KhtER07jm51miQQmQpU3txLXE6gZSqmqucn1SkBlpsIQjDH5ceBwuDO
irrVEE2CPTBkzT1CYxbHZeOvMl+xgict6N7A9c4TAYkTnnybIxhP59jTqie5zbSS
blTUOVgls+EFo3lhwSMbfaNHQ02De+GinWhRYm6It9BHuEPQrQT1cnmLDFmpe29Y
/EQbxzZKlyXfrpj3jnX8wYTMcJymwLE5VemRx+RTmRfRpdwr1tFzNTx5jDi8anOT
g7iDsSeKZETmNCmYPPMx8mzOZhbME9z0cCrAPrAZaDHN4qBkzlqZdg0rijeTZUAn
vEojFj1EYEI30AYObrCLdSI+S4n2AEKEfV3257DAgp/Su7jL8YyEqi1Ak+Tzzj7u
6fWECdS1vMQy+8KKsgIPkQOY1KIAAKWlND+hd6ABq+UYzXpnVUT63wx4AGCmVak4
RekAiBlEN/JUPId7bdvUonvhQPFknLheg2SmF091eYoFWxhVWq4MpB0UaRvpz4s4
ERpT+01HoqjjHaGFkZhBEANYzC/Lzp7wc4gzesCbN/ThKHjyGOuhcMkJj8sRfA41
q0MEsmUJ3mRtY5PAxDBq7j6PUaQi0c6OiCr03anRfDgm23p8mcSd8FVxha1Nd71j
noYfEPow8kCrK/IA6Lp1z/O8Pi+rhjaraSDsaBweU2GdD4XRmH/bb2/YiIPTtMa0
cwVhA0zdSiBYhfXUwFMmsfLFCBIU1UX7jpphge4IrkV+waIlTx5/3PHBSoWEdeLJ
rBQ8UXFuewRoVeY6PlPYD+2ewGS1apNKx/vWMgwpW3cONVn9iB7r16p7W00oh0xJ
kBnbS596FPqPg1OQrsiN4bM+1+RRw2NCR6Wvnw4P9KMxwShyF0OYfPpFBj4dOlTc
BGfOU4gPdEDaDoj69rj4nYVFlnz3UABv4kKvtTWVFr4QbyqaR0XMe6SL8l2tJY1M
FvuVWp/gH1KKnsKa4nSlW/7qjKQ4u4IhC4JA3ve6pfbSee+nl77bDe9abGqEdLw2
vAdLBoJxbFD1r0kAPDD1aQi5KDefiTvclqULzXHe/9D+B11YXVVrE7NnsjtVtN6k
YzhoumxE3vEwxMAJU9OCNbGamYIU9qxVEISjpDyjXmG/Y9Q05VXJWbSJDwTrHwcq
ti5riwnOB+04vLKCzudNeNB5U4eAKOXNxr8xtmcRNvvBHSwRX7+G/EqmkmIdU/l5
TLpCxr21bj3rDHdfPq2NOfpPTjnPuyujyxGN8sHy684AlcxQsHQAOqIwEX9n2yPg
TwCgwQjVmBYv7owWLQsuLUxm9SWop2C4DSAz8/2s7RLMbzoNWWQ7nb/Yd5L0Jil9
zRv5tV83F9ENWqVwwHbuvH+g6uio5RACxKJfLGVqvGDFQSHyeEWOGJtF8wBmRQkF
xaJQ7p36jgMC5xnUSsV3s6BhkoG5s9PlDUQXGqfV9fgKYpQijObsW6XywlUWaUeP
VTNIFD55sL0KvnoYhLnl9AjzyR598zHIOut+D0i0Nq4Sh+F1ocI8f53Mi7X27eUR
DqmyOnJ4yFY/jHMqOjrqQZE8Xh9HxJdAOzvneQG8I9FOPe2BxQQwBKzgsA15cx3s
eigmLRwGG6QWlmF8myaWwpHC4IEW20LdWMQyBmr7lia3rqM83vk1fHYaSB0yIuE8
3iPVYEusF5z+KV/0CTfhcsttmTNUAibGtdzPA2YyEQ8jj2xEQfrSOiNNYR8tGD4c
HDYvBq/GF+npu5Bziy8CTBwDXYGpUPaVu0eg7pbsORR2IfmSaHwS+s9ySihAx/z6
QbDdfBkPW2e0ihRFBWGcoPHNfNmPRZSweLLGnSI+F58xoBfKLfDglj0K6TYNxrRj
B45g1dp4YYNkbRFKoWieiKNdWEZkb1T0yPrTycxfUx2cUIYqNIrrWf8rRLNlSVGP
xEn6YJfh3ByuEVtQ4uo8KgvDp1KPfZMhgE1kqUhnZzUQRigpu36zEi4QFbE76BtV
ixzX1gIBBBctby2pLk6uLvSwOdfXXI+IkcjiqXgWWD4oHJ0GfOtgbdTRpnU9hKH4
j3sczXql1X9Nxfg7RMh6TxkMN8py6psT/SXfemmqOgJOP/SEVxGW/RXYqgjmzrfK
RUGhrl/U3QRdCBIaRH1FRq9JAZqO03h1SfGeY7522bWe+8pCg/IPHeq8rHh3jqnJ
Ytr/ljOetLEpK7zyWq85xb0JsZaEptLqAqo8AKIggz8ouY2IjkyxonHEyvfShJ3G
ldd1UmQldO46PJ1+NIzjsJtHWzVFz5RAogcvy/uQG/U3AeepKGie/ADfeKcVKE0P
+wzfrUl18588CvwOAgd3A9FYtLqw1OVIM/0RA1wU2ea4BYXJKCVLTPEXxagDDIIk
8YKjMx0+ZgcU76UVqexHYrioK5I9cRaOVfPUIXyCrtZtoa/m2d0U0xNzTMW68xDU
WLV3qP2CyDq3f2NdxoVvrLVeuqZGWvzayZZVSHV486OfQ53H4DHQIHOF9KxuGUY1
VRHe/2T+SVr670Zwi5HESBkGw3WLAzzQHBVX4YhicYgHLB3ewt+V8YUsy8kT7MZ6
fnyYKVP0JquSUfEymK5W63RXAb79SxDX1qKyC5DFIwNHMjzQ7KLIHLB1+BIWzguP
dSW8uGabccPSmkXAqzlFTmxDX4jB7HoL9ShX8/Y8EFH9zzsJOO+CCrGNMdixbzw7
JDxEOacd2woZEMXtpkHcvgJfQ/KntTmb5YgjZ+ZghmwJ8+tfqD2faY72YcG6W4YO
NJ2Vijfmw43B/0QHOmuLPBkdHVaVGwYsU8zfDiH/6jaVxUDdjLXZEl7RyG1rhOZk
A/KUR88o9ilGoJq7PqbXZcaSQaSGBrTfnuRaDx6VSP8QlJJukRJ7mYm/Tut1k2YG
oTlxRIcR3jMXqEkQPxrbfpSp7xkCR7pk0QA8iAnxTSpMoIJ8tFksTyVL0kKZrzNS
P7vP/GhihQ7VrE4dZx2QY4daSWCpoRHGxWFF6XDvnNCzYWDon4+YXRNyjT2KUo/o
jd3SQaJhvIkVYd6bGqXHtL9FS0YK+OKn0d9cGskTy2/HfWrvD1rC6eZyNeTgcjsL
oul3aDA9osCX7xsrOi6if0hcqSnb3L/DfQT7fn/zUSuw+TRRoqnoechH+I3DPds6
y2NFxrYpCj3rKsJPEc7QqJ1G+SUy7SA/NLhR2BhPBicJhGjJZXLbsT7pY2ujg5Oq
4EyybHRAHYAlTsyHwRsDuR4eW0QlQmGI3y/4ntubdTevkLEV+jZk6M4SFFV/iNdQ
isS1amSUBAt9JDG5kCbtpMxtAlQ6rjfu6KB7ppWwJlOvW/IJ74QMnlMEfe5vEC3i
DBkY9JJS/Zi11yf5qDE0di7SCH1teGJLNsFBlb7CWrq8WUPedyWXfB7sqr1uT6PR
mu4DEPCCX/oSgZwMSdmJ9qbAOcGuVjhgNpTIp7GkWnsnoKnqWzFsRzga4SEYyTvc
IhIrwyBR34F7k461f/tehYE73h5iLQ/keyGXsiK/yM+PjYZkYZWEU/M1uSYTptXw
7rtKLCXbtGRzug1JbERcp4d/sZndIJ8+QWeEB/2rNfABOISVLssWJc5TtYHhrcvo
kje535AZ8CYChLUoOJ9rUAWbmg/Xu9vxaEReH7y6yk2gNPsgq7wdX0RS6Q0F8Flo
/qcBofzusSGQflIfU9E/1dPRb2QwsTyT8VeUDhptsAeDQO4cy7N6nXfn1hEaU7LP
hKoOVIAgpqJG8znKRQ/FoOgVyM3yuGC2oHy/ZbgHJC0//uwCJsNbScoUOUFhEtTb
xReTznwQFvBCvzNeVaBX//HT7iSk+URf2pvdZbwrWbKKCxsfdGTlWkipdwVMLnf6
HxlPypKg/lD4Zqw5drZPcqTSN7pNhHWeflmEuedfy7C2umLHx0rsfF6e4uRylHMb
USVYGKU+3ZEbhkpG6SIc0ZgEDGdEDAY3i4ydPnDrAaQqmso+veap8l2RXQIoZvvs
f9IgBtyyBWaYM3QocbF8TaJ32MAKgLo0RZ3xtkBfRkzWlIBjir3GVPeyJxkX2OdN
bKzsH+1yVUrGnI3GQV6kV2CRMpFsSAD4h3Jb4D5ZIH5Z2ysno8rZ8Smw0S+i6eDf
/tLAgr0FQV3QXqLVL3l/89VPVzn8AnG83s1ONCk684rmewyo2/mQ42DLle06TjRr
J+4ldv5DcqiIstcCbaLsP4ri+GYKiNA1wT1XTz8V2Jv6nT9RV1TxHuIUcfM9CRUp
lGEGFZbQPXpm9rw0AiPgcngqNVt3FTVxrLfqZuwWe1Vh3gY4w9P2xeuFTJdK2HTQ
IzYEQEMZJSBCQLfGsgEhyoM5gjD59K04e5yaByqXrFTgcYYHFdjwYDaGpEoXT7IA
m+qMxNj6cwg3S5qFc+RPUqRfgnIv4tysYW/HraugQnxH7FeQGpwtJXB5puKgqKBy
1/RkQ/Kki8QOJ55DWrmnKsne5XE/1fhTrKg2AAzhCpdLiToowRrKqJl3Vhz9f8Rp
Ht4V/Bdmczcm8gUpebhRIhLb37hEPY/yfgO+qu0lySZzmAa1itjWEOkqDOywI5eV
6MJegv2nrBPu1RUCmJlbL2d90KIrZRW+hQyaI2/Fb1H5D3OvP02u8Fc2IymFjG6r
ttpIa17bd2EHfpk6YSSqJTLFKojifr3YGjocPz+TEdPrGCa0sxHCsB+RR/vBoUiG
bXJoaj/nIpgQbHPly9oX3xYfhbucpVXiNKNjdJ1JsMWwYJcQTgWYe+da4sD7Urqo
1uwsVH/TRkDCL+oZ4qNsV4DktEVUF9eShg+sM2e18UlYPwJ8SEUwlasy0bICQFwr
w83zuZMAjarTajk53KinId6M9Hy3kzpRfRwj04OjHg7wH3QFNRCNKciaQRgKFQq9
CADkm+os5MYUc7syYK4vp5dnVOI3iO+Af60iGk6WzJVTP497LbUIzFeG/PJPsUsw
NPoDhZLCPI3/L0NvTWyRr3Lzwz3Z3d5O6SEv42yCQr0A67UEaoH1rr+13aCOmBUN
xe4nJdTawzSMKhoeU7qgPLpofw0179bzj7XJ8nKUBBOojjj1OzKn3jzEx3W9AbX7
kVJKzvO8mqtmpnN9+cL3dC9xuQ8f324FCroESQePBDwTrOngZdU4Rr4v5OO/Wm01
qkL5gBaJ+el3mAco57PIKb4jmc2HlxELZlRQpQswSqk72pBOun72pJU+vodFdYVw
U0OSMyvZ1iqxAx/HEiyrJumAiI1Kct/XjGSQCTURDveBNYa1RFshxjfsL9HFzzI8
hSCS6EY1sPdX/faJmvLfXPCcJ53xTksQzHKoOKJcx5d7ZXii0FngBMevo2CwwuIE
a4Q1+6F46E4/Am9VVSnHaAEGRHl64IuWh5wODs7kmCAxlFHfoAdOA6O58eY/3zeS
ReBBEMtwBWjg8df41DcQ2qVBf88zjhSrqHhAAqTAwnaAGOLnC8I4pBlDHtiLk+0z
YUW7/YUd4X/IXLQaZ4ocxLfG3h5GhVikGYGz0UIoKTSDsYWn+AdgJHoyAXktlUQm
Qr/tUQliW9gbRPrHtm/SKieNcHq24qhGt2w7DzCrBBsq7NDbK1RjGglJNxUvLR94
XK6T5u/C2Q8zqGu+4D6MxCTKi59BXqpuQaaLs3qUxG+jrwQDlpU4ITsW/NC1SK+m
aVrGFyfkon4seRNcZiDc6vA2YqL/831hzcmsJMXL1X/+up0esDo7X1dtR6nvdWXh
7pvMYcNT9Fv0SzFka5HuA6jGIBrp839WORL6issh/qsk+1nYBz6yltMvF7mH+WVw
5m7J5uINyZ2xpuFTRNBHjWIsF6+nckJQ8riMpDtKklB7Tf/jTC+GU97GLZvGovBo
YZryc8HOBUqVuJwFFwo6oiEpup55i5zqLcEBsM2XhgDyNClza2QCxS5hF8I4CCr3
WmS9jPSnANTPWYDQEb8UeQ15oDy6CqIoQpHJDQAHWCXU1QLpKYmaOdX8bxKrtRMg
2AuazhNpnEN5yDbRs4lYL2s8SMtlZon13iVfGZBQIQFkvGpwve6/OgoKiqVqmzP4
ZlL5yy+dlrX8UwI/xNj/jODUfBarD4YVMDQVNxte2W3PouOZ9u8gq1TAOjXmYHnN
76c2fmeLqC1+gLlPa+yb8efoozoHQqRdYAQARw5YhTTvOPj+fQseovnbhCByapmb
6EftZ0csJGwwlEgjLn5JImv6EgTmGZziOyC+onPMZY7Z4v43RrXxOtV49VHdCsOW
x6tP1iD+Fcn9czl+uL78WIigrvwvAonHS1WJUyGObun+AxtpFE4YPmo+wc3Ac2jd
L3vHWDleifAFOS3Z9n7jNm6rHtlRsrhrHYh+caIKfyRosxvlJdfAkHjKw8iAUMTm
FQhkGHahttK60YMzCZqtsEG66Yku7/j54jFlDAA22LUMI39vf5QzQIDppRXMvzml
xjQ9wt8vbE8s4kg2d+LMTxjTo9npAtwbdQzRGx2XtT7GA5mgS1w9pK0lNWxP9+t+
0uRV1iNUfoGrynt1nS2NLWyEb2EnIs47pU47ZhhgZCTrevztTlXkptUntojkrQ9Q
WGCeHtqOl+NS9bM3IrONLS2oNXzI4WZiNAXYJ/TTgrEKwMSjQQNwYfu6pvXZ1oyF
MCYVhnVffbfkOki/+ZwMzA/K1+nzzd24mwv/hH4OPc/3lul3qdWurepcm/hH/IYW
EASSTr4cWZi8x0wzQhYdEArNuyOcxvfr1YTaaUb6tz0nCwiFpp8nE8mFW7+W5bsp
K3mUw8vzaF0iGaDujWS5D8AB38xdPOO09NIQoFC5UmDhjIc5V+vJpUKr/RlUbP8s
kDz3dAp9rRCb8S61g7G/07bAKG4rjCM0iBSoDetMsBFUU3JCxdD2kwSPI6jkm1oD
kDyDHS4EO4e1Sv8aw9ZmSPq+hda/Kte/Gl5znICcHULepi0fu75M1i89WE4R+7qq
SOM/W7EOEfaWE5KHiecOdC0+kvalZ6d7/QiHQbSaCmlyQ9IoThI9ntP2aec897U8
JpokY4xgGgjSXxJ74dHVQJ5YeTHipigO962A3KZY9Psje5Vl8G80i9ll0KhHzSv6
3gLny5TMeJHVelq8k+Bx68ieQKhS2YZ497o5P8gMuDVwZKjWVcKwLwrUDknlmU9L
71KZrIGJGjbt/koNNstt1KjfRr0bu+DfAEiDtaJGVXzgbzImeiqAZ3XWtE29pZY5
R+IBHUkFLE8sen4TdLcp7xE1HBvwpD7Wa1WUoUqUlEM0W5cYUGnjCYQDEfoYQ8MF
gWq+PVwCnzsFjHG97hrYHqbK3G7UUAJrYuyrbSoW/YVukB/tujhy5kxac/QSzBgu
IPOocUg5Vtunv6TzjNM881bVpQBLZ6fTn6JGbJ6HYK+JpM93HE6ZRZkecb7TERsD
Fl1U5mdiGTflS0a9Lh6OWaKOKcl7Sxs/btLjy4BAIOv+zcHoYb7m0C3JT4RpLZ5i
ykoPUrYbAavCR0s+9tZOEYX0ntnecux4wApkEoBS8ZSntnJAW3tdKFY2HLZV1tsO
yGVaB3AWrbNxdC8IlD2T5dtW3vthMzLINBD386+EsgZZhv/Q5we9YqxYQhtcn9AA
2A7GQpmaZEtDokIQvY0fH0QQ+MAvZhFcaXIcYMnEey8lWVYV94ZwrP70XTz3bpC0
ysp9x3DVbGdJe7NBNngDE6+5j9D6S00JOn47f7Zh5JZ87WUosbubZDg6wCoOVMdi
UWfvGu6revPq+x6P7H/M3cHYbYZX8V9IO/8kKcDUbqYBwjIaHNGBn+vpw9/xAG1a
o1m10/oLsMqx0KBoxw/sRxGVfLcJzQ93kG7RpWJCft3d7GYe9argkVlRN0BhoUHZ
MWIcsq8pKoqj9ZPw9+Dkw5T53yrnYAXXh5ZLHtU44+5rf8mMYmg+vXuGf25anBHr
k8Dj5VpiglDBY8wVScL3iCQNlnP4XI6Zjtw7AsG/BOoZ5KI/gojJdYWDVeFinszm
133j+krK5Ivr2FraULbO2j5fW14M9azZKtCNKiWNOQ1j9fYv8s6qKsBFvzGeEs/g
Y/13bB/yPjNaytpJuP5Ji/BCL8abCdwzv+EOPOSXlptgR3QpamKdcZ2C+uxv8zVk
w4qbpiowXbspx9g8NIXtSwHIfRlmCWXFUyQCEFCk1PA93fOv1yKMkSy2ND6v0TH/
ZhXRSBq+WFN7RXSWWiOTxkUieaqzQwdR/sc1eSqQXmxqgensm9NQfI0idlmM+6CO
fO7h68p6esRWw0unYs8dfjnkO14dnaLAaugtIIso+A3cWNskjshnBmzVPQwY2nL6
Eej6rcZLJLMmWX6ehDsjA+BApK+Dk+fN8iz6vvESLMeJg4IlcYfZTn658ZT0g+aQ
0CgZOTwxlv4VY2YJ7gmaHSY0ZaG0OdKb4rxbJm4/wiBxr8sTiq0+yKmiPCsqlGDd
3lbBE3yCYZOPH9LobwlhVxoJxAdCZxaiU8R2+Y3dvarm3vgymK6mN3JhRj4NOnMH
sPcpZunfp/21m7iUM05RvkfnGu0yKEuJ8r+mJfdebdBF/mTsSNConM7licoSM48U
/2ALCjrawP8Rf7TsOk4hbKthnDX27NkkIxBJwdCabg1L6TBtx2HBVeegwC3C3TeB
jjZf9kacoDPXbPn5/R7quzQe2bOT3AwkdW6Vxe8LGVQurnU354sHbQ3HLGG9MCds
mzNNMiMzgc47uhf06vikAig9C9NCq1RXERBwwhEIn38qRkbtE6lXLYIwbcuPqCn7
iHxrw9Ay/aejeN71gIEGrXU+QDKMZ6wFJ1y3DVnbm2ZTyjXHnQjX9LmYVlmdsH/h
r2LQNLDu+ek0pVv+hB5qZFUGKLy4IlwH3UZHPzaVnHzVZXJkCPwHm2VvnHQcDnjf
CGx0dapim/ps7EsI6z4cb3SGgZEg11fP9IshgJAPQCY+yNJ9Jraa0eaj17YlTU4J
bjIAOaA9aLMRZ+1nrcL9b6hagDWbjeQZvxOEiXBPeIRm5ZR/MJAXUPPhPS5VMWaJ
MIBjVHJZ8E0qBiXFg+jR9Otqm38kt47y3IT1M5ItgbiT0AIB+ftvuo6J3dRxH4yZ
/nIDvRIEzud9l1Z8Qywv9ZQeKty2dZ6B2XcYBVRFrrPHLbeabtr+B0ObMGFP0Xce
e58pRKHqReUM8czbA3S2VG0O3LSOVgvX8ZVpS9oUY9SVowr7YwiSy60XZ6KgAiGf
tvhif5G5uZXoI95xa/uihOyKIt8sSfKyEHN8DrX/3s+2dcBa36X1cgraRkruzwoQ
PaacouhEBCogC1nDTbcZHELvklfykPXByqWBtscs6B1GsgP/77BDnVWGu4trBVlf
aK7Vz2Ptfc3kfCSOt0CDuImaHEv3gIFuZLKhrERxp6Lw1F8E5va01mOZNTOcaRp0
HzgFnwz01M+h8t3TGdusxYvqkneVJLlxHlmQo2czlPYcN9Tc4BtFyvKb+KD7i+7L
5w9BAZKP7OjMnf5x0FQ51jrCvOqFecZ7GZ6FJiIWdOdQVapk3X8rflhOfDlv01v3
GYtfUHMnYQgdVKLPNEsmstxKzrYz+cuv5e4LCf6889+0w+10stFCl4u1qR7u7CMW
xQi0K3AVx66bF91UZA8I0V+wK8p85b5ZuhX7nxaY66zdNhcR7aXsrFSZMGkPQETP
sqfRGEHslmayrS9CnvZtGi7w78VCgcLcFIrCKTil2pa0JduQoE8A9VeQ/EtABIes
+JOnYpZyl4JRvOnoN/QIJFrEkO1qBgsh6LM9dEczsGYAo05BtdUYK+6JoZWUHrMb
FIcGFoknZt2ufX9vnuNLY+RO5pndPxTwl/NEi5xdIXddW8Xn9ArJTTh34EFrdNUx
ejqVM+vj9bvnk1dKPOjdiQKNVbZziPBTdFQVtigm6lsVgB+H4ywZ5h5K5f16LjFO
m6Cyz+TZ73DuE2iQFsIPSIZVCzuuAxFWkeudjhwmweA7htHbKgqA4j46S+EjyVN/
+uaAZKvMfvVwlxCwXIROxC4ElJXAOSgdWSAGqGMLzn9dshsWXG4Czkb+jukZU6cp
PIly1iuQoZNOjUg9JEJddHbLzJC4Q3EMgMfrpIm3+tTohqla9PnjvDDZvadwKlpm
n1rPu2F6XY4Sb+QsqS5C0g6uPDXSgUNCeCSX1KnbD7vmPCofIlf3AqLEK6PJas2Y
9vl4nfD0IE5ZaJRhO3fZ6fMVTSJvMpraOYvhM46MCsAcOs2rMfhFl7gbzePeA7sj
6YsyzH56PceIziharuANcT5gwzp6Anu5fhQNHNBDAZxYUHI+Niomni7/noRy9Iau
SIikzIlwYk0RZZw204JEHmFQaeMsVMH1q7MSAlyyol26kb54lNLDJVZ0jpgs8bHW
8iifyKvx1QripSlzULdkfZdlBR8ER/T+XxCCAaQvvoM+9RYaQd5eWy0YDIZJ/oiC
PxtBqGxQh5lMiY/GhXrayCe7nn6j6f9WOsZwhmzwHTbuXWCMn+Dz+IwZeYngXomd
1R9BeXUT8G6+pYRV5L60gmassVv4kgpNlbfqEvWyDPt+S8kNpN9LJTamlZWBcDmF
ofLRILZwOSn2TXKC+P2U9I97DWUndr87ybD/O07r0v0OpmTzJEqx0b7FKMzDOYvf
jw6OG+ennv2CG0E4XtFgiPB7Pw6Z/BH5wWTvo0p26CI29QGjQSt4633l6YwSMe4v
UBtV9bw+wAyecd0BonUs/EX4egsPVZtOcR7okt/1pxxXjZnumFqV/HQXalGUH0Z4
rAKiOwAtrWkl7KlXwnvNbZRzgQMXKXAgqwAAge49MoLFGGgpR7v5X7AWQO9jPScG
oq7boRSNCSuijJniFa2qmuCHpVFtEJK2bYVs0eQVRISR5K8u/TUNlDqZbN4qKpAY
1TPIbhjdhHAawVubJpEXEo0Imouabuv26uMNglv1svDPg2CxhHkQi2P/15ipLPx8
jREh3XvI1zEUh1gBKLBUa2ZVTAdMH6Pr4ahZJxZJidaXEubLGczHNDniq0SXtGxp
+9j/S9OckaFLH3bOYuunBG05bxP6dwQk29x1tq65+i6d7z5xoACQY8HIquqvFkmk
NBYtROf4MspvJkam4aQbadxmhwSfNPbRM8DtZOS+a5E2Lhq/eBmBdA/f9/Q8EFCT
kfwNwAllLbXGnQFujAhi2aNlXRo0NZvgvGQ2OrQISAVxqkU7nzHcCfI48tshcDRq
qubaT0+kQbbmMhTa+Wi8cBoQ9NQhnLTzsoegJZ0RMrPlXOt1fsTpgLNihW34/AKG
8XBzTkBiUJrtAEisLe9GH4T+dTK4sFM2rNZaY3GeDDB9yT8AeqgDl+7gpGpzqDTc
HG55bH389q6AgSjE0hvkIDYJUWour38gCHB4VQClMkfktSCHoCvI7faYqwAvNjqY
0l9kHahw+uidPqpB5ay5G0tZd52X2RajG5+nBIXfrAr+6W4PNyC+zwr+8aBk5qmz
5/PbCe0pMl/0XYofIfA4lZWn/9JtsKC267SxV+AZW5x9CK2DdIH46A92xCyp2url
QY6Bw61HuGgaWgYLR1EmpzjnU3uYASbokblbjiqdsP2SS/v2awPV8Z9Y7KRWGEa8
3smadVRL0K4JKMQIyrZ4bXt/aTkK7MdF3qfwMkyyuyjayk4/KoxDOJGj/rZPS2jw
smn0BOYUZna0aRJ+BmCQ5N3pFxA6Fr8r0gD+KWOml4llzfK43SsW302EeMLVgScS
87iIzu0qVl6PzR7Jb54douYwV2r0ZLgm+nXmOEjGfN7kNB5t84oG4evqqPsl+XOC
k7XJ6o6D008S3znC/7gm4dS/KOMXa+Rr35n34CrBpqeKJrGBXQID3cIscKvdqfEq
a3A7NG2REzBq9nmTchdpiL6zc0Kc40kAh4J/1uXNf8bi3uMRvA8Cw/SUrjO47FNN
IcbnDnjcBAzcRQp3tETPLlt61Y0dKm1GxCZcDnp/okPrxrsfVL2hIOD1P1uKuYhK
bNgsy2yzMb2gOA5EH+YKDzeUlexoIrImQNDD2XnYKErM3g1mjFo2WJ8AjgxcpPwH
QksMNLjBwZEeOUvZEyzr+z6Wm4E3lhK9dRFGv0TeEG3nuoFf7K4lCxhhvYKsU5Os
79SAm0eB4hO6mZAtGuJU24S6mBmar4wo51Ym2p7OZ5KnyepMfh9x9xtXVomSyBCo
YYhXbcxejHHDsub7s/DVqTDO/K8zeNrh5ZKQEOk+DzTOVShb01NO4RSQaVUI26Ll
5wVWhi4R0Bpn6Ssw7w8RoYSLPAo9wfCNitROk5eGn2lU4b9+uMgV7rLQnitmKLe8
dW9WZF+OvmjbOzlzpLy7tQgfaYRp6xPM65ahUHeDmZ8nFME8eU9VPLffguKcTDTy
4LO30ZfxUQSzk9/x9i8i7R9uxFutjJQ0DUPqowqvCKeofE+0r7zdLQIPXvr1yAzQ
EYr37pKx3d8tBrYGiryuX0TnDQKbMa+0sIerQhgMBonpLBBJLxJATp7oztO7fQta
xVE6WQszw/EYyMvPTclrwbThtuf8g+ZIexFwrX/TGPJBhvOeeYhxnEMblLI1LQaX
M8vOFp9MN5v2mqeOpm8rtpSZSfF6YWEfuNsj3AedcycB+yGNWmNpRWEI7CpzOnwG
VFJeHcVROkjCuBE0oTtAd2qU1xVo00WhxVNtND8DhNlAtbx1f7pH/qZtVs5EV23B
RqNthmoEJL/I4LBqrishwQ7Jc5O2BjXmSwWmYkmrv3d/DOq2/W30sJSeqP1e1rHx
SIp+aw48QzL0ayBzEVWJvVyq9NqMgSSwOiC0lQiVrW28fAzzgwNl3EOVAYAKr+g4
XojLOblcnmVI2YzFnWwj8nmqZB5EMNB+2R66nQ3ylEkNZVjV6FFI+eP52Z1se2D0
FAxEYoSq6grqkrH/mrbG8DU38/kXVA4WInS9UZVTB8VJgPxFp2hF9oWaqixHTKxF
SH46gY5X0DKMvkCBJMl9R+25HHeca4lH83BuKUiwzL7gcXgD8vYHa5I4cfKmZ4vW
MA9SYERjp7lBewvRZKL0WkJzVnx8gkKhT4N1H34N9l1C86wOT84LxYvCMCF4B5dU
ILOFaWwW6dVPUt78R1HMlFmcN8k2CI96+ju31u/AKVw3bpiY2itoTAZr6GJPgIRL
hfIuN+otPUrPV+o4FatTvGApE1htnI8qWTWhz6jknUOi7JpTC+iR8R2IQNKmGwUs
bIXMuUKYn9QHHlmMczCjrE7Vsn42dpZMSH8Ak2Hn/b3kdLY2+nW+3oMrX6lvF0NY
KSEDo7xdm397asl3rqtg1Qi36YxSgLogN+JcquJH7om8IXJWz6Cz8WY4Q5HJg6pb
L79MSpB6UrHQlNGededY/+68yUnQsuNWoosbvTbf/RJFaXN2Y/ejj1bTgnxcteOf
/ZuS/p0bW8mUQ76lZtIybNykG37gZNxqB3kPGJpY1sub/DbIdbHR/4kidnLR0cZS
2/toAqHH9lp4jtamTNkdcsOPNcIpV7q6UAKrg5FgMSWHdSKic9BOBC86wu0/9e/O
+auz1UhgpKNjxsL4CV1FuC571mxSKORzdb1bzmnEiewOwiF932Jz+UEuwXf3sISj
MDz6vYWopQK/QNjxS0dXlkdyJWyGZyHYVVysiAVvbrgThjW6NiG2QWL9urUvwohX
8wqYSf1Zb3EAynULpYH25zkaVNPHKjX01n4K7ObOb6FN/8dTe9KFfgN3dg0RpWdz
81v819/ZONWSTEGEabGg29M5OINyUcf1Pe80JC0k6o/0hGDK6ypyuHPFUz/uMJxu
ho5pVVjpcF3dWZnOKg0yeWhfbUbmi1PnGOPgyMhikMQfp2q4UYLRWx+KBgDUTPFy
zi/Q1LK2nT1eRCooatwCUg6hf1MFl+wrSCSWLvLlg2FGKv/w5D8joHYFQhmpDiZX
NtRC1bgehFdfkHrqOyIAQWG3+UqfzMpU7PxPcDD7KX2bNsDaqlh37g+Z2ORwgUWY
bmJIIEdMct7IMr484wMCuhueX2DPg9XfqcwKBth8PN64aXQNaNEBJEzWeZR4jmHy
1O7FwZdkJ3UFNRxrFvHBJ9FlFGiV2G8wE6vihMbgqqKWJ9qXKYQJV3LgcaonYdgJ
wEM6qJFkEZQ+fNEmne8iGBK6iA/mvRXmShVn9tWJ1FrKkCeqGWme5EXQ9jB5nA1O
5y/0jQx/XhngIT0fFjRYvHGfU5rih2ZsE24sv4+zUAigW0pDJMG+AjAgLaDEaC5b
7kX1S/Hgw9Ox7rRjYXgT4111MrPVwRFCoZKQYtxewvCccMqsO3bdZALAJRQdIJYs
EgfWZef7q5Neharc3L47He9hpWYhf5ArlbMkXNZeVSS3Apd8KNzU70woIt3YBoZt
lBrn4zPrnc9eR8szp1UbxBkvQlHjZq6+KvIQ88NN+jMTB5aqXIgLHfBV753Rc5tm
HTxAH/vPhw9dqFsGSZIngjbpWROTgAufcJeviW7eMVS8Wapsvu33zhH32qs0xJhd
9N1IXxlyf5xBW1gW0NYtaeWBOZitAC3SNuwKD519nRT66OoMtwzymTM6UOOe2XYc
6NHyZUCdOWBUNs5iFnknOm6k+pkPPT4GiZm6lFnjXyK+D1rDE6WJZl9j9uAcSgTj
ZsS+wFmhuMWFOtrNcKL5QuhVZPQFFLX+iUPYx/oOOigzN2EzI5eeknQiK2kZ3h/N
ky0ip+/EZJKGf7xXmb3s6f4mTK1y3VpMMho8qvXfHGoP6kxKgcYKkhxoLDWHit+C
0p7dCoxPsGP1KiKBfpn+mFrp7dN7noRz5ojCaSxs84Dp9bPLeoVPc2p4WMM7sRaX
vR69efhkhAS7wRlSLqcvIrzhUbjLoA9e3b2nAXokCwG7tp/8Wthi3XNJbg2C3nO8
zepEDCr2BGnrMHTO+d+G/7eIC6bj6iMtAk/dOFzxR49e4jiJVJyvP0jITWGjB2Yz
JNP6hM7Io+KrTdzGfx5Izuu6BGVrqC0mAKTWfdQ2d3oRsXUdnHIipUCJ3EdOWMNM
yXgBP7vY7ImKiPLgYRz7y8t9MKxte9PJ6cOOp/M2AA6qF10yy9s6agKSCPVQJLB/
lgol9sektGEp6CNwWm0deU6DxYwie7W8/R4/r0TJsSpz1G0iLGNY3b693+hXIlPL
YewmdVHcQFGmFRt0Fq1EKiKI1JIyiUc/hlzwVWFvJJ+g4Y+McoNOQoFj7Rqm1okU
0OQxMxKMy2DecyVpf9S89byPe2sne/QWqoBNVpsVadSNo9QJ/j/1W80yJBGMPG9x
KjZD7sXOD3uYeXT6z8OK4HLR8NXpog8+TqoJaBcH7XrAeM7c48Z1JEWrVHEjm9Kx
1jj/iDk9SMkyRN2+lEK4n+otfOL5EkEAXN4fpLZTtTDFGrZNwrNmXyT1E5CGFub4
h+6d7lysCMoNgLIjTvL0aHcftdFJB0Dmla+i42BDgNog2hvIjnb7klb9wrUi+D5C
61lhy2ngXZqeVTa0k2WmL0qsYKnrqTD2Oa8lxk50z2o7QrXHVvaf1noW0h+AkJkx
6Zk/7SY7dTn8AIy1dg4vi+8IdcrN01mH+hh/DHO9Myp9oxeZoxWk/KlqvkBl83i4
CuVYwc85jFa9qQlfUiYuejzvMk9IBZK6plF5cNJxVCnkL/l+mCkqRXqgyU5tf/hX
SB80BJfzu6+cI5iUhtQEegUGrqIke4CSOZfQZi0JUTEUzFuuWD1IuV6PRfFAMYcD
XsqMbCuJztFI0VSUOqQKuzXP5bawT5nUGm+kOzGIl0jcFmOb09yL1Uu48gMjZWb4
hNgdwRV4uS3IiKutRAL/iyUw3YIAvkcECPV3uZ67e/eUM+GELMmE84IhY3JaMS6y
T2rqrHPHJYgdQ1b+pxrknMuBxQXGDroI1E0vc5CW8bWozVJxaBjywMx7wZStCYbu
bjS9sDfcJaZZTBtnStzOZAoJQX2AxYSgnWrZU3MMnjWeHq/S+bXSP38i3qfPg9wN
048m1AGJc37nq9uvctpgF5IjSzQkqsPehYzFWdAmKNRNlW3FAjmK/D0oTsqBWAKr
Q1h1pxHl0hVHSNSvoG0OphqwCQ3KjWjLwMbmwZ+o1GLhtHrrMKpJXzsK5h8UiVm+
B+S/emWA0+ye58EKGPEx9hMCHHOkx/C6wtQIwQIIJqKs95L2UYe5ayrlYhmQoEMv
p8sgFc9dmyywNgbh6Z6Xe95jrzouStikt0nH2RRc0bhGjRAF7aUyL4jfJax5FwGO
q1Dd8y/Zo0Swif4zT/ncnjQ8ohUemA2qF8u33ZKHK7sFddbbG4VbqZwQMVxLZBv4
y8Rii6auH3c1d/vX/J2wlU6crv3Nj0JO34acCSnmfIEKrq+OKMNV3qTAYteL8hH8
jFTWEE2DRSJhoN2Z9VEoxj8UfLQlidfJwFsKbOx/YrV2n+UR1ATUJcziBcZF5RCv
qaOJJ/GgL+WNSSD1OsctnqcRWMMDzgenRLVAGvgz2LxvosgnjF53A8Hu8jN+dU0c
0f1KCe8ABdlOs3HGwcPU2lZWcYT87aVJKr3LQC7nGtUu24qn6UGZM4tQO2b9uO4C
ufd1Lh4h9cO/xmjTyY2kEvOJNDSgkmBSxw3sCVa1EnVtBAhnniy5jxZXSEiL7N2+
Sywd570T3CO1iJ3LYRUA1iXjOqBxvT52n09W2XFo4gM5b8AOTckH1BdH8Kf1QTRf
kpzIKUvzR7ysf9/V6H1EKdt3ELpawMMO66AB7JTuEsMdIGoqEVgos7csXmlAtoFd
6Z/BBsi0dfolw5qwrw5pvOHs1FF8xhFC5gWjPRqSjer9wzPLSd6LwMdMFsF7EJOn
rF8CjeORuHd203RKk1N81io1E2oVTVzoiYeqKb0Ee7AhBEjt8hok/VQJiPulP4VC
7WjtGLiNF67dyGBUMZRYLxWJ8trU4FZGc5AAaaK/kyi/dj3BdMb/sKBfcV7NkoRd
sccQ9dMHFe/+pWrn+NKuPEx0SK4ewdv9Bvw42KytUPGuUDjdNKR2v9fOIPhmonC+
VECCMSeazJSmXR0BeO7AGCxxOdJ5UHfma/BRV0hRMsYq7yqIozjs5YsV/YEGCm1N
rKTYFsUZKUXHvKv2fyPmSHeVPePWnaa/1Cc3eOTYX2FFhG9I1rVJboD27MjKT8nz
d0qin16hxAG2Sy3Cq/aA5IZ6JAhX1ErXX6ZN5MkDwS3ONdrwwMTmmWJahAcqD8Pa
G3gu4l1QUZ0Fw5hrLmvVAw0RdTzXmO5gzzOFZNiMkEVFP1tWXwZvzmfSpUA+QNl9
g+g/j5+nUEIEV+M1Dx2QVYDptvE7NP1BrJzEiEmIOZvjcqFDQzK5adZTDq/HzVqL
nhjAr5iQhiiC7InbqdQHkh0TaWRo7rjc0Kf+Ra2A4w9dLP+38kMnq3Pd51y0wLjc
TTtK1b7fMD0CyadsAW25zfVp8a3c64RXSyIleAUmLiWcTgOLug+ZayMPieNEVjp9
hVflMT1vGHXsnBLtEP77ON437JKK6pomOjECYNB7+/wDtocsCJ0qcsaL9oUPS3C7
64KECVdKkfZdwgh98fqRle34pxeslyPes0gWdcf7Kj6RtG4LM4JiF2dbBdfgNjBA
iIjnw20zMILgpc3u0iNhjCIgprMVJQ04whLTLjSt5/C/cy+GkDBKHtAlKzvOH9OP
+1PPg7uCc0ctL+SdjcASOB8YUOG3OypOGcl+xAhWQEkNQpbjqO6F2EukrjT0EYLq
5w50kBNgRqu8XcBWad6Zr2f+i9nJEf7qPWKcMoJN4Y0L2CiypLktaCz/PF0m42HW
HIdaHy1AbpHTM/YwigVPv31liHAkfGe4tPieFUn1NFxKYUDRC+t0zFbm2sL3TwGb
eQYKTSW5AZdjx3rOOl9bxwSVzB/PO/SXrH1SeR0h/GjuVKR71BgoZz6qWGVobo5S
bcT65ljrWPpdjCDHIkEILGtB97+nzsWyjO/9uBN2knNWumb6f3q2dLSHGpASJySe
9+cKRW+g9Y1hTEZ4gY3Ww2Udztp7MYuNPzTZvh+RDbYWVV8VF96+LVKUW/kdCKxu
5O0tp1LfwzTGxiYjZnjPt/1/MvBFuuJUSAPJ66t+dpiZQRykp9pB977gwFOP4d+8
hgs+IUVP/lte+PggN9rhVJpysg4pZVFNpWq4LxZFF1f/H667xTyM7kzCN9uvNAiU
8cHe8X85bEuGkQ8NE+svW1p9QQBudVmKr0dxIFD5ur0euYzgW2zD3hBk+qvpG+qX
gu6PM36Bhh+Z//cFxj4igAnyrY17QJDs8yKn5wSVCjb3leu0g6GkFP/ZBxjhosKy
kZRWI0FS1StkcblcCnNftF/JvjEFN8XOjPpGwqCEbchMskaLmTPMeFJ6LRPcNeac
1XMSlfDitXMEU6tS1TnIEJugk11h0+maMiFixC6vYbKnUKCtZ05AnEN3/q4GwHIe
61uRUfxFv/g/C/bsP9/OAHWEVDRCtXLMgsUMyTL+GKJ00X0ivq/Q0aXBbgXjBiPC
NqDQ2FMTtWJg6GqIk9+brmnroaZFc2w3i0avpWmBWk9+JBtachEu6sY70SRvsWyn
bruRlUk0MEFGh7ez5zDSbGKdBnKEph8TlbHdPy5OY/1uwUhoCc5/1lD5cSHuoxJp
SweN5wCr6aj4w20bjGRVGPUd/hPdn5eF8ZPMr0JBE5LnaHVTewT7nyyDg9xIaLAb
AqM9x7h5rvLcdo/hRhhWcOQqwvNbnoFV4qLHNRi9j7gos2xGx124zlC3mxMVupdb
4MRw5oRjBtq7LnI5WTgiKoZOMUdEQeMONG6TuGk6AT397kRnjIFN4xK5V7OSVAkz
+bgPuMiyNjW2P/uVAOTi3fGD/K2iks+8gG5DZyCZjamzGIpaOjTPz9/kG6NLlrcZ
iusz+G4uqvGKk1T/N3Ea5LyxTNTdxWjuPIdXRJug83DnrfGCFko3aELi3Z1W0Pl+
694w93dEg5OLZhedMOvG3e2oOAeWPJxnFhN8dTYBuuqJrjRXkaLf6NEET4qZW4T1
FFoEcH75C9g8vHpHlZ7k6VfdXJ5gDcP2j1yiKE3kDQeOfRv6JyZxyqW+COvu7O4E
FTA9swqaCHJEsB2dILSSQbJ+S8mrRSl6i52NSPck0pEsi15LJxShCjxZtHz6107s
xL+uws94bgO8f6ztsL+owXW9ik8TBuIQ2UUPXgjNTTPv03cUlAJ6IXHnfzFPMXd/
kRvlKyTkhNgpElF6SE9cIlQpIURNrhwsjvc+i5IlCSss3nikpxC+pyOKuTKJ1hec
NBQlWiMubKWq8J82LX4dfTjBvV49nMpUspHURVerIM33553zwjieGcfdPbYhGwBh
9z7R9AruQAGvgJypEUSK/6u/B+hJOJblseI9OzuifYoaq5sPlprOxb8Tyzx7GoWS
Hg+kmMlA2SHKN/sB0CKRgoKmNMjG3QviIkmrHKj+/r9g+DueTYAqFwVYaS9OIzZp
2r7imBu/RASiw+tYv4Ws77wdTKdNXIFYA/icb9d21WJ91+JOxaUOrvIcU97oaUBB
duP4jlrAAi1wvJrVh553MBPJnIYAVYMGVOS3cg1XTWs5tn9y609wqGTOj7JTdiuH
bGT0tV4tHczHcnn4kLl2ECHq+vjivkSId99u/wJGXZFN3uPdCaiE7qpgfd7hBq5x
cMJIDYlbjIEqAO2lbO7hUQf6bQYAK8dXlFIrTdDj4r5OfhlmSJFGYw20iWadXgXF
MYB1X+WY/M4pl4ppi/FegdMBlDt0i2X52WxgpowfcX6a18GSzDjcXvBIiDbV+naP
FPTvOmUts1UejdFQR8WcNtwxiogNhFLdTN7L8TALpGabNMk99VQHfQ9mKgUkGFCW
wefxW6nQC+CziBFF3nsWzh0ywurfZiHaYbuL/3zd3F5Hb3fCeTxwOzY4NgIOqXFw
/ijopcgdCZhEN67i3KXXCboewKGQExxzdgCHH6JHvKNR0vML+EXyYVRR5BZt3SZz
8L4u7kgVn9RjVBWf9gf7dp4mzpsvbUACzwqHWpCraPLMdweAhpMHZ9gtN84llKSM
NCqs0r3ARWndEBNd8kX3RMHGST6E9MSpRafDW5GI9K5CiF8N32Fijum7ntvNS4ug
TflbXbJIJ9r2/7ZL289ucSpw04pdSqGgF5iNwexsQQ5P/x94m7lsfVQwzj+Fjvr1
uWMmRtQvLrhZm7AIW4OLCH1m9S2fKsyvWYHtVn7lg6roydopRmP1xX1sTxKhZwVn
7C3ePWVeV8c6GVKH5B1qJ0UDCU34JDSxkUfcrx6noqUYr0JMPcBNqX8swVz4tu6o
X4i9IJDEdHQHSZjFTtWnU4QQU25+0xEMqGHECIU/F+DTlrEBtz9RXwTV6iqwP6yi
N5DlXD9k+nbRvKmJQRqY/XyvoiS8f+e83vSe4p/GS7K7k6Ubmfp5tMqPXNVME0de
S4se126mm6Ubz8X97jbomH0Ua03Lcp6JseI1VkvySsfxOvHTjjvXBXOT5bcO1GyT
RN1t3ceYr34SQDmjl2Q2CEcrIIzeCxAcVO7RlfAmq9RCzBPaWfWSwdKKppA+lshL
RGGIOYhY3gdVAgLZ64aeCcJhVqXjO/sbwRT44s1G5owPAtoZOKLFgZxTeU59U3ad
TrRywL4MIYfZtfPOV2udgMnIjAVTuv+IsWqUNZVnij2IhM2pHHFt9g+suhH6yuBA
Jc1k7E6f0GVgNcAL7+4WoNWwngI3FY4yHWxME9+mXwEA/iLo8W/0lgRjh4WP6Uq1
Gen17chIpr21OrvGWfb/gWS+mw6ULLsQbHwAdmnTu3Xrkuex+VYKl+PF/djivtaB
cc5zm1h9KzcO1gHnNJZofojfcH8iJmIsK4xRKOIAI4bXww5S/7CsT6ZAaA3PHrr5
HOcmmK45yHCO6M6Eoz6OCZIC367tr1Zv5jIlGUpH5eydk68DA+49isOyDQYuUMm1
FIoiNt3N2m1XKcFZyZlkbURcLsBLQkzqZ+3Bbqh4gCDvHAIoJC1ybWBHQ0vptz1T
xw+rkT/rejyTCinGA6TPfsWyx+fZ+v7kGlf5ypq1UmgtD52X37cnWocrjgqcd5M3
S1BBnbW6MH+tNkxRfejbvckxPMs848OBlSGGSWHHnUukshDTuhxpLAl3UfBfitrL
whHgWlCrzuJocsZBnGN82pHoh0FQy5jI/EngVJXvmNVqxkaVgpaS5v759amhOThC
tWAldup3GOZVPwyspVTllhHY0zxwAZNMBsyNkcTP3RghPspM0Gkxx6JHYMOKN2Xu
sk+x/SIdJ/5tUjBgACWhHYbHJ5EpLnezzBR6fIFAfG6z7tesyv4CyHYHXlqxt8JD
fRR08QFOFR/9A+Trv3Kg0f1gC7JlhxpAWhfSTMv4IOpPNFXUUTb95D/2BI6HPeNM
HmEzvDwyq4D9hJcDqTneJFVRSjHVonvlq/lKAl+CXwi/tpWvQWVnIwcBwCMhim3R
2hmY+Lg4B6kdR+XDFTkiEluewyqu7jop59insJt9UNHg9yiN6V8tYqxkusMV/X0q
LAeWOhUE2WdXQTGzaGWid5ipugHRYCtnIGXSEZWJktc4eul4VxwqTOntJGjtIxmq
1OkYJnlglhh6FY3rgiwg2cCk1Zqxhhfb10Z5vmgTEt+4q0SrAO+STKbybiOg3ZEd
+V+sGYFE6yRLwz04fyQkMD8zrHhLq7uFPBdpZpNqTqNlbgbNyunweeDSQ2nsiDZ5
6xVOftCTKjfJYmlDy5hGOmLersheBx4goCzOUfHwjN2GmBYWnnxCi+KawOAjbNPh
COfyHWjGEKH4wakHeW1DxbGHcNsqzqI4dcP/zLGSEDdzF/jMvBT+hmTDSakBrnVn
aQcxoXrge/d110bd5ug540IcSRb6ZM0rYiEBG4Lv6Q8paAyaIjmwQjvHMlErwwGh
jkp8SUKZaJ4CSt+1DjcjZrF87VKr6XB58ujRJYRv5IvuPueMTU4ZGkdseU+4xP73
wYYTya3NPyMZOqvhY6JdKl1GvAUaG/wNQAhkniLgJvxind5/QSH6ya8xKonZVP2X
DAv7z9EQt6A8GcMeZcZw7fPJOxHzXFEuotXWrYBzDC5VfHSSIUhZL+iUq1EKfXzL
NT1i6pUoAJi5/n7ZwWoC4bQgZJ0Si6Soz9vYLGh/rY5ev/NoJ06foE/BH373mo93
+tz1TBYdmvqzk+WSWnXRAgOCbN4dVXaa7iKb2/Z4OAA/g+NSQBa1tbg2F813YszW
fZNvCRNUp3/VLG0jjNlrxfPIC7xhQ7EgbfVKk+EAbG5/IXmP0mFp5nzytXR3g4D+
faf01Z36wH77MDtmQIdjNMoVok/qxkLWCaAw83DeyOZuhsO6+YKej+diXiRHAYur
KIpDS/3bb3DYmZdrzD+wkO9XF91BPTrIhP9ioPOyPZ/OoJbgKPEBI4c27ufpimXi
Ovja/LqRbJbTa8tA+Fgkj4NUnbvEMz7BmSYHJOHqoGsVgA3xhlkocYRlok9dpity
aV/3GNU3Yr4IVfI5kChLjXJByXxnohGGm4tP6cuOfvtWrGIDzZUsSS5cVkicF/NL
MgigxEzQC+ya9Wws0e3m++eUKmQSbeEqCYsyWFN+9qgBqLJae8UdnFAllJ18CBtL
nSrCjtJzoTg20ODBKLdAZiJzpchtIvjy/gVqs7Rm6V7JiW7mmBeQU2/MeLLVQR8i
blbrrW5/e+nfJZWRRv9A/3956M/wC+0VtMOdl5ystSjZJ+B4B7AuRl7XzWtB0suQ
9db+ucBwhmdPRn2GeCiXqM0ZWzrFbkQeC++Ah+4U++/rG6fNldbUk4NaCcjniklM
/tJ14O6L19U28lEIQ5t957lsYUcvHEkyfI54elxziD5kc2GSdxlYHzzRVGC+9kpu
8buxtuAssrQsHssP1nsthDruDacr+rvHcDqzggsXl+1JrYzefRfr8PEHkZ+3SVAK
EeDfzd/4wJ7xLTbGSbMpN+YGzaUBsdKS3eluxmWt7REnCeOC6BvUDROCjNctRd4y
O5dzULv2TaEUPYlwD1I87GqeGDjrpfksV/lxZntqLTzY2tfLOKt0BqNla7//sl2Z
CELxwFTnWFBUkb80BAY0Y+/nd4mxzIc93qoRTQD3B+ngni1REqzzA6ghP1LLGDNN
OlQIwRqwWGm6ofP7wzAuRsCChM5Ag8nodmGr0oR7N3iB/7l0hcK0s8EDriLIogI4
4EI7UqcdrBDBDxYayrjIdrFNtE00WAaBysRW8BHPxrMPdutZs7q5L2awJF1QtYGR
VXX1Z/UCXuR26TFUcwZyFBeYuuWZm1Pds4a2X47ZlKy0S41j6B8pYTvTwqPo/aBl
iAPdUVIHvoVwfha/R+dW9C/N+gIBGw+qWV9JhqMnZM7J2B+GegQWL/IrajShVOku
8T0SSr6cUtb0wbGf9nLQN09tNoqhJD52Wth9+UQGdU2kS/o+O1UfdrF4gSGj5kK2
wjbRsWFXRuTe7E12RZwv/plAOceemZVkrjUoPLrERc9yKaeDKb0sVyGLbNX8P63a
g2J4ENI3pN6rks4D0rZJxgaiLnBp5CT3qpetrWfWu8/YYeTnc9PNK6QyPfLBssm0
zOQEOKrFNyNkKYWG6WXM69n2QeuiWQdtBfBo37hDvbSN4U4awXbr5FuBPbzzOlwO
SlRKeJiqZfOzosYeFaDs7cs/rgF2rgkGZJPz73iRO2qe/6VJweAa1xOVGPotBaGR
6v+4gHsf7cOiY2rdKjopN022yWEBn8oF+YJHmH7tdY7erlMfZGUN+H4T89ODhU0Z
HgOqAsHoM5N+GQdj4CGNrqOM+Fsri1dOEMAfq73msBn/l38VPprYswSmHcLTNqF3
LslXGEwtxq4HopElZgqvBzCbEQfRd0LwD3VnsC01LbjwXEDQj/2rcOwnKMh6cGZl
pR/aAbMq5RliUJSYcIKylBXUlrhs0Ym19RC6TCud2fB3oHhTNwbIcXWoLD+YlU7N
EIS+ymqnqpJiq/jigGGpCFShUEq83Pm1Fasd8eb1/4IQFjfpAOLmyT7tAiQkfDmm
zka+QAVIeoCexbPL7qwxNOuaynszxbTX+57GEr7fXBCBoHW+sgz2ed3IkknNoT6x
eWz10XHUEnthf97Hu1SULB/ps0tHdGASA3rR/MSLFfwH/H+6PVtMnNcNvAIYlVD8
M+6hwQ4RXG/6O1/2zclfFRnNC5VtRThsMewEcOGmLodzQLUOPTb7Eh3+TkFCjHvR
so7KGXj9h7MxgsqdljrZU04Uy3F8Y/h2t2uaWDAuMZ4vef4rk0QjQA0AWpBjmWUE
OmDgPde9YTKbNZYSVGwP6Lj3CTI/QQQZ6D8UXFyNpQGLlny7hi3DfvFszScTX2rE
g6gwnAht1v0HXIhl//PYbFJp0eAKMWXl1c94i8S61MXntZx5s1d1zXX10/dI0yqc
m9RzesH8mo55Fn4l3ba1b+N6qWwsoSIa6yIkByd1d3CxPtIJz1HrKWiypHjMz02h
yGbXze9VykjtLWg1HmZclQBtzKvME8cOFVoaVdR+R6l0QgzZFDBsypkitudx/9Qt
BNyEicx1dfSCLhg2Xf+pe4GfY0dInpvb91fqvyXjfGKSK80Z0iynjBKL+A6hdtE8
tmz09/MTe3yPby1iyt/SrVKAQf6Bp1JP6AEpYw32KWxlQQL2UWEK/fmti+o3iJwI
kdu8MZvFDWC6G/3pZ+pqNBcqEwJnodNaz+pbjh5B8yGhWDeZw195+EyfEQrIwrjZ
dx79ujiu3LbBBXZ/iNn26sSURClxp7PcMx4RsKn6t92J2N7oVYtw3buywGqI6YRj
+tIRZo8ij+Dw4TUGVD2Np22LnKbnurAC3Io3frCVtVdspkdXKco2Hwms/gWWy3sZ
lv4oECzHmhA4i0iyWQE+5u+AUy83lU9XX1hgt2rnZarjYZiL8DmU6G+1ANO447Xu
NgwzNuPmdhlQNzC4J6Tlm/IxqZjZs0j9744zzKuMvXnuchn6Ps7ORFVa9eTy4pkL
KANfcr+oXOa96955zW2O34ly+VGX+JKl2D8tc6dJukQdEkPOJjOoNiHSfkqX3yvk
8ha8vimnkA5Iyw+Ff35PfNmr/L64lXEOciZaC1wcz1hli0nI02ctPCXhLWXM9DHC
X1McL8Q/aOBFH4CStSD40xkdZSXQz/A/KeBpScmeKjC930RdP3N16cvhO2G3RII8
PyHwILe1dHhmreqi9Nqjz9cL6hQN6T6P753iKhX65xaPY6H4KWkA25uXN8VZnYNx
RR+2mrQVXebsEz72lQ0sBceYAVzvTzjJBwDvWXEgHGvkBaiuZI3WF60oxoYflOIq
y/BHb/mw3miSW+1rkRQMtLcmB5h2/qlBNXKpV3gPbz2MKv4JnhqA7SQUKtTkrKMA
2z1hs+jCL+oZrhDE8J4unFxrw8pmutjtgkcMO1oKtS0CCjOjE3xeUmITo610iB3E
o5F3JnmOAdzvAQl4AnEnOUBuiNFHkS5C6UoS4q0/eDqor9CEICZBEm7sMAJ/dyu7
0xI3/goZDP5nOjM2q2a7Vh7bTSvcYRei3DCZP1uxR+SOGk1juPI7+ZhoF1g4e+Ml
Jk94mqZG90DP6EVjHohCi+JQ/dNoNVIS7mmjRsPDID5twmj842uUgSaba0AgDsyX
ibmA+b0rF/ZM9zOtH99Wuu/jnt7KuSudkCZEsO7zRF1mFUEnsbG7njF52P3ILS83
xwdGK0DhSDTA4IRbVBddJWHJGHGGev9IVpvi+RDaQNI45R+9cLh3JUImJi7it5qK
2e330HgadnrZ2kVH3hvWxCaBrEw57OK+ysmEM+Pfb8x24U2k1zrHVUIBS7zUMAlY
ddedm1jPUWofUo5+ftFM+z/p60n3Z+GmLkTzcp3/xH28bKrGWUdSucTwjlPQaJjD
CZpW0dh0kHZvyFTJQ742xN+G5iLAm3/qnzCKyGn0uqXzulUeDnYTXBhGGytqN3wB
dL4H1EIi43grB09YfunPwd6P+Xue1NMmWVbgWwxi+T+GgD/MAMCKWd6TpMrAuJef
2rO8GC0gCbBP1A14H+8amzQqPV2s+vy37+WkDc1ugPVqvRzb1OTV+8mc4NmmBXUe
xfYUjA9SX+/g0I+3EzkfKipX0CpQwhow75nyzyyp09sa7UvXoE0Yn4+rYKYtdkkg
xkmIUHF4UD4i+ZtxYx6MrfB7tTo5RkMxTaph6S98Qg+8YtsCk4Vco5Q3ZOBWWewu
oRfd76Dw1u19iYQeXcoD/cY5qtaknLF0KFEzwWwhvlhdvLsm9+XLK3sNOIdmZwzK
sYSK2jyOMijrzvl6zbU4S/2TkTjqfXfWgruZsxULccNwnM4h3H5GWI83Y0Ax9b5f
Nj2nwPIhuzxDcp2OtutJlym6fYg/k9s24rDQsg/PQoP7DzYvY/HWr1wcF7tM0+sj
9cnKAIhdusCc8CoKPh/NSqpm8id3dxjAxKOdAHmhaCVdx5Q6ro+VRjzEtfoFR4ma
zqVmN4Eu4ayhRefPyplXT8eC8HHhsNOv6PFMDWWG5NF7dJ9Iv7YMYorccfAjv+PJ
+c4vqVFkFGNQb3nZBbuRUaZN77it5BfpKRA3TpmaZ4uXZWnC2qkb6dY1TWvTggYS
RpU/Crgk7QYinMjaL9ST2nQboj38OE+QCPelHjax4V69EUFVLNBCoM8IEoXaxZA3
euAqJ2n3FZ4iqVxZ9hxjeoBzeYO4s2PDlIf7V6gnvoSRjrOCIrbvXwPEB23HKykJ
iJaTBzh2zmE2pecVtRuz6j9cDdTEL/iPYno/L3W+2K3ea4FoGGV+pUWLH71S3EHH
3p5k/ZvSDcAXH3DsXt4w/xGwRigSlrlC2oESOnuyXNSD5//TnzUWF3TbCIsjQ8RF
MkYvTpjH5mrU8gvWN6ciJuz/hDk9vbIKVmGwZghIzGA0Ekk9tNWNCHKuxPuhyLi5
e0Ry4XFmfWDu6KFH2Xqa4g1yHFSuuhdPi8hqKRV2fHS9BHspC2i2y86kHX/6SQy5
jgCNpEUveOB28l0cyicQMMGsVYLOiUJEPSRSygBYrOLBrZ3ANhNAUuf84YNB4Vwd
PL3Xy+XNOv1YdGONIZw6X086HLHBxkwHVxNHbK8GRbET897RXB85aufvn2ltiF0p
qJp9DK73BtzsReEbNeVWFbcz8OpDbgRRujCOj4/pqFvXUq7xADxxTZAIvug9JT02
1R3+sOwJG64GNg00jD81XHJGT0FUHbaopUA1U39Mas5D7QWjDnYlkg/W0U4gdB5U
TSdYHwtT05e1M/A76BhxP7oXreiXgDDXy2WYwPmPrxXyefB7z8dLzFiGKZku9VSU
nifdwQS/t7ykvqvdcHpelkTevA2PMv10rQm7bus2cR0w84ImYVi4kSPI8eTXAYiL
KXo2fVMFfqY8R4P140WYvbfdSHi2BYzZ1LeIGXqPec2BcYxCIAMhsM9VafbOw8Mj
1SKr3TAknBLsBfvn0m6CCQqUbEd6n43HyRqQTHzx9G5MJXuCKak2wor68j7G2Fua
suepy/xAzEgu7OW7FASlhFBxHpPce4KYtgMOrr7FsE5xEm0Ir4dbvAwwgfrgN36L
exBVGyowqg0FIQVUYt6Nh8HnQjX8nD49HaVMPsuOiTDl2t726DKkYpyNudBUbfRx
Xra2DhtWQroWAvq99mjIhcxZBZyCu4AOQ3cO6oKoDLloRP34FOlQwuvPj3Hme7Zh
IMBM8vkslgIavFO0/NzZfic7c80pPFBql3nWa6FEPoMNC0gVWAl+MsSk6C0wb0To
elgHHhUaFq9W+UXr2ZWPOHBer+/usWYOduGgCa+kB+1/XiRY9BJnFlnGpaeI/V7n
7+0YMD+gluDyFmpgrtUlk1vSO3RoYpTl42iUXEvXVBAOgjMp15AN+9fp+HJYf7ES
5o6zungRXFKEZa8BLXxW6b3/urERhngSCIUu7SjnYKyDO1GFvm7YYA7lyf4l9P1J
0NT7+hDU1LRDzMQ7D7LEturralb3CWsa9xVm0dfr5lCo4buD9+wgYieDOyXuwPiM
jPbmxUBgV58Z89T899wjahcd1W7GtuhZTbPRKo8upNEXBnZhb3GehmXpfVO/A2nU
NG5E//S3MkTEYjD9+Jj8LU4XN5QzdW+r3VaBJaUa0X/tNyrhKKuTankl8JagIl7V
2fJcD2uBAEjTvgHIXLC46GxliZEG9T2iKEqT97vQlmm6Xsn2BvdyBaJBvDH7uC6o
Z7rllttwgqnf7HXCsQQqIJOJum5jI7sBpasqtPyX/a4/COG9P2veFTcZkLyTCRgO
JtcPfvoXD7EuCFevWDuu788mlvyGGjj59szkdmxZmjYjuARa5J90T/dlhdhGIMXh
KTubnyH/Ss40khJiruai9WGCD3bByK/zSSZzDtk18qNp9EGPFQ1SmwUBxxAHOdu3
KjHbwK2dT6zexrMf5n5dOXZdig/Tx2uM1KCsUX+j/ovJqvZTRH7S4zZGX/bAyOSe
lP9bTiFqfeyX9CE4BBXsjnt2kVNqt5jd5SJBnA0kAnlagDggk2lZTSGsCvNdRmU2
BhliC3qb+h7trxlg5elby4JrswfGg5xstgRdvfeLjPsjsl69JgdzSDiDFAmIEd1I
IkbIyeq3Ik1VVZunONXZhsVZB2HZKvfOspVgFCRlmrM1CxbNAeYoh0YpROIxUopp
NvvF/gmPmx8YfJ6ibtdOQIbCfcVDkEz0QjNuu8gPo7xtUCfYfqdnQBCt/VLFMQHr
OutiVRFagFG84h664hBxqaMIFfTwjDcn6UWm+pLBr/lWTuz2wVLLo9LnTLCyyaNi
+5SG99kJ2vgXjmlH9RRiUzgufu4z1BmBlbhfxR98W5kPdlApcnpdC3sUeUY83rfW
uVTZum3c+aGkcSemzdpmf4ZKvMfb3TavV4Muoizcq2X7wc3MbOD0DPTvFu4YFYfH
t8ccyABajfAho4s5CNFxFz/w+LymnImox1lVe0v2JjDkbZtS5aVxW72IccQyk/RS
Ab0Vbxuh/ScvM825ydNa+HMkj8P0rclthisyhRTqz9vs3DpwM9YoA0ZggFnWPe8O
hkNZCkZ/fWo3m5aKkLfQHSjEFjypi3o3ioLFbYtO5anBOmhTeu0s81K764By/z+S
Hum4L7lQbWWIT+khhqzl1ZmdTi72x7DTKT1/uubRc8T54gPxuRygiTvO2HM9NS2W
eO5v+ped6aHQCkzdW4nQPicfkzRuvTdneWEvTzmT+bEiZL6AtRjJrX2UhKwWHWRP
b/I5kVUw7/ZlKNeCiicddMW6r+R8tEPsX+naJlCbhNPjSl9wRTWX/CEk0bBvnEJh
2oZ7tcRyW9zD/hAJa53mbrnciRTo/57pdYQKv7dPY1zEfrhtvQj/+tHAHPZEBxmb
NpvIlyHfR0HLD4+g1x+hGqMLdbEs5kubcjiMtUzBHUXfsvrJyqOKYzplfaAVQT0D
PfSFT4IMF6gS0dqhknEmx8VM30gFUf0ScvCZw4ohaB0NeD5XkykO6HnEC7MhoQjJ
SB8Cvf2g/fQJ9VebLDVHM194U7rZ5bW/HFzRtfNytFekkCuMW4VT+MyfSBszeT3d
BsxN0rX0RjrwLh/tXIysN8XhzG3Pc8EsN49kfme0FgN34zBRjv48BJJ8ckuhpaOg
BAUQsqHQFZYiHJMZ+CbblBRdx34fogzH5pEHeAAYvO3SAcqsMhQbAjDgBLem1kPW
PEe3Rx6G4XVtwov6wRtcldILnfIWqlK8Ecpa/7qvFfOIjOjPTShFuKIAEguswvlQ
l8lkvfWjghrjlxmOyUxxNKcNguwyilv/8T+WvMpbmnwCsk4kVN4CuwHfs8GqMRPV
PK1yCuk5U0OuFz2i5taqZb+ANIBhG5ln9ToQZF8QUyTFZ/G4JaB55C+81RfIucKD
8jPLfdX4G2PNH5rOeQHMbhV7w3iGJ4/E6hLTuUpmEBAh9VhvNqm8P8gUntw2ZuIC
TeJMi0Xr1BYbN4xe8qP6PteblRel+nTuHXdBbXfeRkJGjXTblNe370kTW8iHtIPP
rKA/ExpQNOxRR9K+tw84GVt4EqALKIdojJb8+TbxuKQLt1zGxgC6B1DJgh0Aw/gN
seT+7kCFIKCHK1aZZonP4sR7weJ5Z0pnPI1XrMAeN7wTjj98ZUy74jUlH+w+1+Iz
dZhpvA0PcYGndd2YtcZQWQuWVFtskHlQw7eUgjF4EO0/MQPWxsr2chUkvPRDcuAV
FR5m4adXAxn+WQYX3FKoeuZf3oczv6AqjD8salF3A3bRAqSmxtHOStf3tSSf+9Dp
eqAtYV81yRNXTAW4x0QHEJyBu/1o0/0ToLSQFeV0qOerqWwCIxkSt69RLtNpUenG
1a3D0Ri10TB9P0o6NimDCC4i2hJASsyy4lmCzRoEfFb6V+rv2FWcmwTDQHtN9mr5
2EiG15nzmwC/2CZH5kUKN39hX95qKUPORTeTOx3UatyQIcqKR/+gsvRl6aiXYGZd
l2/dk+QE4VmEglQkzI8Ld3zLPgV+9p88k0mOTJKrb2d9MRwPiFkF9g6HYhCWFhnd
4cjr35U1F8qJmHZpnS6eNCzYc+3Og+TOwJkB+dkZ4e8de7u8kzQDiIpy2P2NB+ex
oMhbYiiDJcP+bdxExgozJNlV62Brjh+vhmSb1hXvtZfLoa6mA5Hh1sJwkQKchF7E
0xdcZkC8olMCim3WSxAAgugnWiJvpNRva8d2/mZItsHZZX4tPInw4G7gwF/xKmjK
zHvzQUXprQ0UVaEnxEfBfyFZh8KUDHdkITa7OULcVX21BMQq1UZKDUuL7+laB2MZ
7X6NLpHjTO0bopx5wbYsuX2Lt+VEpymObE0Rj5mILbwxO5icqYrxBQozEq1warQ9
sH9Tw2NBoA9FgpX9Nn9fr0wIsyySpb/LBy4ET/FW7Z8F3njYs684Se1nwA3TteWR
s8/vXy1TP/Y27Gh8XaSr6KZL29wOVzkEK1qIfXDa1ugQuIn3p3HhieopS3QMy4kN
ThjnqxFQChCgQNHCER+px0NcDGOjg8hGqwjsLl+dgGDx2RAPRZExXTmm7cadifK1
umCs+42lfK2Rr/CP8J53lagt0lP+qFGSLjuP5WjHEx/JS9XtKGsYza8EAh/TjtXK
I1dC4ikhZwu+4CYoom//6zYQVL6gyr11gJqrx274Wenjyu7KuPhXgPvkfHPuSgZu
WHn3MQbY8f/N+EKwC7//ZZr6S7Z4e+LU6WO30Fg4LkOXbC8z56faduPdbtaZxaY9
e/hr1NzoUc7rTmAQ/waL8o5vRl/HvjoBqAlXh1PEh6NAWr/bCjORrDV0QZku+zVp
5vSZ0E9I5ztaqY8l0s3VTKjPZJkr9v3HIiUb0z4+fXNsOx15OzqjrNOlL4bH/Ab3
lz8kKJXGgDuIB4iT3Y3BeMyeXcTRhtlBgpFpT0OSTeBGZdrXdeu5xkPBq5tHy4y1
WBgOPmQBmGV9C8sX7TZf1Xrr9cGk0cAJsFgHZHLPSOYPXj2azpvYZ8YXiKUb3NG1
N0jzlc4+bFYuZw+41Zam5TNJZXn+4SFvqBc3qxYfn3FGj2rWG96c9OdFzncHgxIA
q/Ww0HWkOHIscfAPdDMHP7CNrt3VQ1waEKjcfCizPMtLiyACdrekwZqPnCJsAJ0f
99frGjLDyyW6zmoaoUHR5tzD4vZCXiyXbZ2IZ8g4/9gJ3nblLeRRiBKO9MXfzp8k
wLaWgu+98LOxRUlZDLZX8cCYLU5/eAp2bp2SyWje42Ptoh5L/Wyd83psfY2EIDph
Fyz4px2ck3KZ+keCSLaA6h0sGU0ES9GH/Sg5FGIP052mbdb81raQOAstDRW1p+c5
oVowFbTVQRnDIlrEuZD+N5J2tcxe2JLCGepo4LLG5RgD2IEE84SQYfr5p8XHu4cK
yOTcEmfdeYu+0IdnLCb6r0jeHBZQ3RrEJtUZEHNiaQeWANOuT1w8NQTrEsB6eSc+
jQFYKm5dQxhRO/5xBm0T4CdG4ahbNlp/n4GHpuFZLEZHnnRBCOwxm7ZQ7cxwMLzl
fRMj97jgoiHHrDhdUBRumkCOJyMyePF5BYLhDqTqPc8wZ1SNkEc4sZRye3E0z/lr
4lA3pVFVs3tVFP7ZviFN1HDjZKbiX3oOlmUloH3XVdksuZhneTBCs8vjPGmf5xZK
7nE3/j1uCVZFMUicIHz6QcDa4BPAgSkvqX/emmIPTkRW4zOZefYO40p6JxaKUhFN
cRYYFWjKsQLlIzL7PX25WneFPY3V9pmuKpEL2pVwpsgHzUXaaplYjTObXLfiSBPZ
MMnsJS9BXXou6JFoila0GKwCiUxr0VWG9g4haHwSMhlKJ1WPUlsBW5Y7Ejo/BW05
4Iw9EcMqb3/qQJhZWH/EijxXi51tcdapVcq2wL1X8OcU6qtJDDtflY7BzXlmJGSn
KXrtyWHa6GET2xpoPUV/pWEQ7vCJ6Q9fOAgNSzaW2Nd0m4kZ1Ttj1AHexbGMAACZ
fI842koNDADjeCkSV+HPrWYDmg2qL22c+adnd8ssbx3U4YQX0QADJGTtm6TYcxNy
NlK9XVEbJJE/Tcp7soXvjj3XoobUeTISpADWUv9SjCOZkjtAom//ZQBtA/m37J1Y
1Ol4JascuVtTVTXjRr+wD5qf48px0PflbZQvwrY/fDhcv/mgdyBO/kugnLuotJXc
U28NRi8S5/nUZVJANY810r6WbeIQHTTkJ+vRebaEATQ+iwyE952T/byYynLoUuB8
NHxF1IpPvC+ouBi33vOVG1ETif8U64PLRSoy4L+zZFX/aksqnNRuYWedu2/czuST
zBDATNGGrIrepSfN/0gpjPykRVk961VmPFPeA5l3UpOn5K5SZklzuel3Di9UUdHK
Q7sTVSs+colbIsfxQZaBXWcrN4Fvx9MK73KifgoXbZrWA6AaIbDK1YybEYiJF1rD
BsHsYNpKIDRA5nCTxc5qkPDDpYyGspnRZG0LWaUCoDe24BRkjjRTY7Oh2rEP1/4o
a6DYuuieMD8hgK0n1SVBwhoybL5/Fpd6FqDBKwR+Cp+6asyJ6fa0ukmZKj3nh+ZF
DhhxZEzdBsxF1BXq2eOxv99HBYXRBv7Deg9o38ABdw1kdlhr572SDDvb6iEvN0/x
N5ZGA9Mjpms40m1q776gyj6I7yqxoexnCIrpTaJjY6hli1XNoz/1R7pdoP6k3yl5
I4ZnMg9EODj0UnoeUs2IjxJzXTlYSDyS3BQFU/C7XoSjySry2grVoNP5gq7WjznC
stKAq6wyLcXW1zLsy7uueit8/NM0HyA+Vk4Jyje3fPgP2Li6mMPzSo7xPeO6ou7w
77sVZ/VekBFGkrcrNLOR2+o21fAb3aHWQLDyzWKS6RYxmqmDQjB4OIWaUJlLb2oi
Cb1X06yw0o4+GyIWxoN6IvyKR5SaZPmmOzDEHNZLDsQlOBHb5qegC1b1EwclaIsj
8u86qH2LIK5DfgmCPhUf5X4Rs0QV6PV8DfeLN57lU93pran7tdRjptMcecCnAg66
6udppJNpQEmMEp5icxCLmwQ2//1c2uHamedR6LnAp6iRxC7CJZd/R1m/j65++XLL
aZC67TPBvHtLQsQ/9Eg4a/30xICK9JsYADFk5Ibyf46viXGDiFKPcOOTGh/nLclz
oKfHm4TbwpcS4qVeLZF9nJP9Ka9dD2tBaE37mDeAvAcS0Wehd8yqines6IpYGu4R
RF1VomrDStZQYPI5hli86Ua4y8vuZ31XEitABIVeVYxVgQRWHZ2OQoO8k7CHBzD1
1z2WzIiGJDzDskHCiSlqQJCk+yLS8Bpximv2khm1kG8bpyOwBAkdTihLL7LPDdmR
Q3FPA/JP7WBjT5G6lcUvX6MSEd1TJSllc9vcD3uwDlmjMFW5ra5ghgRwTRtp9MUQ
tnl0AOkSZtrveHodTEo0Eyw5C3xQGXDt+xQKWRz7YfpfsPvTXbWXo5qUGf7zncx2
Ih5MfN0F+s3LKNq1xbtPh+Ha4PYFvl0S8FMvWKw4CxN510oC7Xebmw8nMywZBlLk
pfCSHdlFJHYmszifgdXebX1lRVtMLKbV7NR5lKIeS5mZ1mHIU5FTNvTFK3lKnLhP
luwRO8VvNsmyxDJjbypDI3OcUEOlcGNCTNVGZl7teew11kTbZIuPzG1pi7zhGpa8
RWP92XzufuR3q921rINoCKUJQHfKo7051Cx9HoWDE6rgbCny7o50PllQmyA6g3uB
K67Zjycn2D6eFkRYTRSIpcIzqAUiGE9y1RTgf3eoUcBK00SfjYlgE+2f/Lja4epd
ABNXd9dHfaGpGtLk/hzFCuBW9h5OsyR+gAfr/SH3Eiau3c1M663v+FHC8hGX9K/J
EPUZRsELldjnXcs4Iu0gQ9XFMZZ2XVwBpVoqlk63ZobFzF63BVZ/xvxzKuC83ysV
sH+cOC/E79r/hRbiYyWXACzz2povSfolu3nWh8WBTiyGmjzAzAyLL06zA8kqspIH
J1AIzNoJwesAgb3NUVz02iY06KAsBDtTVkSIOscbjpUtQCc5jjQEoLHAoYFOYy0i
MQKo6yqQ2n+YpDgYyKqQD9JmvyFW/sxMudNyMB9+og/XUlTvBA1lAVWZgCwla+ry
7bcLn6zLljx8Vouki+awZ392mkFsi5UPECDLDMshfgxaPbFuWEzMWclpHcvox9cZ
+ZGCaYHtyhby90f1AgxaJBp61hSDsKz4h6eZeksIE9PlWcaP4+z3RQAKmwl8AVMX
CVPMG3w+NJQbRD3VgWh9mxH5YWemQdNBqb6tnhVUqmZ9hplLq6+9Kz9rkSMldp0R
VddPdDKuECRllztuiaIhiNDz2fxVX/VFHAqqxMux/T0H7LxpIwEpr92vOsvZ/AHu
3Ew+E2R9UvdN0unu8ndoG5QhjCAFZBVu8rZSBw/z99kFcuPvTCTaHMKixl6CRYik
DgRE0QdpMw/e2dNiR9IxLkLDHLnvCADGU6LwaYE13JFVFECc4p27rK1xIlMUSYBj
0HsDJOmGY7jj9AJjH1V/7yZenOnpjKbl37dkyMbh2PDo5BOhREdvi22A0q83nHkT
mzLRdN+3EOdT+hI1cBmSyeE5NdJh+UWuCrNcaAhFLZ6TW3DIT0RPoB8blZGneiVT
UxxSUppsKm92HJlZGMrCb7f4QcOcslIV8ZVlyAoCDzMdSG22jSOxfeafV2TKn9O/
NL51iYXJFch9HrPexyZoE/s+gZyWIE0UpEgc9guUrxYt7LDi/ebt9fap9eAMQod3
RzF+pG7GpAEfB/Kp5n+nk6ZuAcHlenTYEqAqvS9RGS/g9sPugKSncGdwzoK0L54A
BpvOIZpEu0jtL6q9o7eME5jnTyy7GbP5LnVhcaCYcsoV7l9nxlNGmjaCqRkx05LS
ztxLpa08w/5CjJUmMRrvlmFdolxrPbIg50F6FVcMC7iVA1oKWMq9yjGchpa5cDAu
4jkzDNMUQAOVZK+XyTuCfJ05H85zeCiAAeM4Se5304GJtMwrHk5iAwND14cRqlcU
AilsXJgI0nghEbaPp4P9J0JlCmxM5QRRrk7iLw0n/Y1WAhNlM29mfJKb+/ab0MQK
fLE3Ix598i9yIlSRB1vkptuIUMa9UrEdJAL95kyckWl3SKRw0wT6uBMyo9Hyec6L
aghvBe1SjVOpuZNbKt9o1DQuCqPYfBWrtV354c+3NRTJLVZcmGobCJzDd1P71Wv6
VooDWkRiX7AIBkt9U2QvUBVHfMUveGcAl/yTeLbuvcfxXV8JDSIchtwPXmja8KgU
XEL/kJOivuYglOjuF7GPQsHwTWkac2kmfNVBP+B679xtpTRfQmsVGsTKuAEoBDDy
UIpPdAzUh+xadA7MbV8vqixMvHDPtTTzMvgt/3Qw2viEuWyzg/slR/rCLqFiZv8V
c73kuMo4ae8wAbqRjxFPMmeY0CXm/zl51Dj7JzZbIXlvmgAat58BeUMLCum+TbSd
De8+nZxKaY8TIh3bBzaBFWArzM7KWu53GNG9uORhXujTCp7++K8t7ZUb3j6A7UfN
hacLNwRAmkYMA9+SCNd07qUdVPr0S0CMrKyoYcxiWo17dMlxSkqYTJ0GGUl32zaE
HPlPZytTSdjcSl77EB4IPxW8n8nkaNgUHLwgkajHCURAhHqJYb/dVTtngap1uOHM
O/uppaVzB3/vMp9d13VEew7p6nqgJCdquLrgU1HC3YVsGnxIJyi6G91815EGg+mq
C8fGYtAGxP58EN3aDn6FvXB9t7VG8Idn6MF0MdH6DsVkfpgwqxU202nGjV8Rs79M
bjzGqKNkZ2HFSlTEhpipEmz7aYWuq4eq3/eXjVNuEVwtUrX9Jm8hF70657mduhXt
CAcKCZb/iNGc8bCUvrKDBTFCH5R3zJks0v9im+0BpIYkGFw409Bs1E7GUeu7yPD6
CuOde0S/9Ijnw0IidEh1Xrkk75GjX5Y9WHu+OKquFj9giUwWI3tYBcZTYBNQTMcT
kEgSl3GjTm8tjzfHx/4SfOE7tFWYWMrX6plBA7VoAVfj/OQwrIcJ/qNNgO04v0Z5
fw7F+FNjsPWIV3tZMYED+dT18dOuXeOExmckLJ2K0LXqSMviPLVMkix8lYx9YmMU
L3vfNwjY6JdJFxawZBECgXJFGzWtx5eE01NpKJaWx16bYrqdREuU14kxej0SYdZ9
XmHM747MV1xRyb3KoksYyghU7zw3B2WXTpbmMXV6YU5U8tj6pizYs24s7nZrnU4+
Gj7PHS6HYDlHxL1u2YPB+qW7Nj+wUVmbL0mhE2L3HgQm4AQytCRqz+yJK50qvUGO
gy56HscPeBeW+vmKNS1Z3La7medGjjn0L0e20KNWZBR+VTm/96FLT/+PI9aaaDRk
bq324pX3Lns1psItVa9CgnFDmOkN6HiVEJLpiFIluumTnkTrZjSxuOSGjmjQJBCX
UbowVFi6jfTOp6XxSu85KuuOVzlP/9d3gSALd+G9HhlZ0UhmduRHaiTPxtVD0fI2
gOXczr2k70omuV+a+L5K90xs75/9U5xNcAKSHZXMUf6x02tNh0H4lp2HrynVQvaO
EI3UtMaAolXWRC+C9I8wdKHm8bITklJCIgaETdEmDnjRLr5+6ZgPFtpuQwWitBS7
J4VhFQOkjSot3sOmuLUcswWYvv0kJHvflTuzDoxudSBqcLrfR+eW4iNi1FJGK56b
zenzFvq9YqQbO9chFvVFtT50pLZPvvjeM6enyV+aP7RCdiGNbcssp8+7/rJjOkim
QQO6ClXC/uC+nHlr1Ew+0Uqo8alDWdaejfsv31VzMc4KpuCiD/EgrSgYBdIr55QO
+tWTS2TyFYFgNnXxjoUODs7dbvqjKPOdDRwxl3gweWyud4vT2XsjhhYwHXkaSUDS
9gF520BeFMSrCffpJ0h5YEg4IQqM6eukrsjD9LWiq4qiijPcDvHAdlc8zVX8shhY
uN233jDARin0F7aXY3QMZVOxLukZD33J6SyTvRU3MBc4flKmXpd84oxynP2GwdeY
dnpXekRbuV5jwBu5woVfKqHcNIwdUUDJqCDzsVMs7k52lbrVMuwFbvxDVbIduJ8T
Vi9M3HmlgNsDbyKTwq5jGXt7lZ4sOSTr16Er40t5ACxJmLTaHogdBfbbxIa32O6j
LoP5uWSkrzSPlVGVuCUzAmtuR1QohIgCudy/OcFS9btCircvO/N1QCkEyX+N4Np8
rmfaqLJwAt/dlp1T24rI8zzCDzyryHV2E2TtsD2iqHrhZY2u2lXBVRkCmEVM26xk
Tqlc7D+ABiC4649ao0WWxQUvBJZnjlDzAV+kn0Mz9RiMF4aLi9sJCN6HFtzKjjqX
r3h35FEXCtK6yyScycvpJI4rlVaMXDbau103bfzWPg72rfbRmtxWJogzBnzyP7Je
41MGa0xKOb+8kvHJD4om5GKrdTrEIx92Nf1DYeV101HoWPNHPkV1AswZE1T8N/4E
MsdC6iQkn/cG5g/V20uU6HqpIMgkMYq2ZJW/MMZCllvpehzGoUGZqv+Dv2wGmASd
vZglCaVBR/W/020LEbRSKHPmXpJWsQGuQsNsoDLhFxlBab+kQQQTbDnRZm+yPEvN
G3w+kMw9iBbIu1+N9NszLf0EH8RWJggtgFSycAyrTmqt4U+heCZUylAQTsSIi9+L
aZOB8TahZGpBXaFOmGZ29e9TgaRewm+9kdV89lggdMZ+euYaTHl3AdyAoLAzxF+d
rZ4ihH6uS4RG/IxbfXvZdAn3fC+TS5YBFqdWEOQ7CIpDB53KpL1AEQnLuaCZ9+S2
WNfvKbPOS62aBp4qSMgJs/Rhon+vnECD+qv9BTvZ0U333GurKpF9eIJfqkVJlr3a
GmPo5z/HPzsFjXUSaCWuyau3TeyVQg4S4nRpYw9LFY462aB+Bi4+GMnspprGAEtx
YxAIoDbRPcyD/2ggUTOQyz6S/7vmZlpZR5R/YfPM/tL4Z/6n1TyW9n4F2rdeeomH
V+95f5xQTzo+CayJbyhq1dXhpVjsGBx5LbJ9CgTk7KG2d7QXKoIui8xsPu3kOZpb
hWWd4vxB/eE3tvEBqt3gY+Gl+0NgB3f3uLYNNwx85lYjvoUJ95mwmfHDD8vYYQ2D
1lvuOyn7EncsHSmfsH6bkNbmGohoj7kUWD/rsN/MNC+/G5PAApfZp8meq67EfV7b
Pgjiar9ArpKPHwHN+eQPr/pP/eIlMPKX5QXwQ74hIlEylI3D5pZvCaRUPhUA0+YK
ryhm4pTW0KTZdGWO6lARGVM6b6wpZf/x1SoXGYU5gyGtDAcV/fmTNBqCSCIPLe1v
Ojy98Ip6WdwaNdBd09ACYbHzSJ1io8icNveVYetTEfPzz70mHLKyzjkm4AczW9nY
RlR15pIvHrkLjHXhZ1iZ6YlME4EKM+5W6OXwwCXuOVRWtg73px8lU85HdlupYsd1
dZ8p524LGkx6qyDyCQ98KUfOVZJ6EJQgrqE+g1pKsq7MEiSjQsJowjkuSmBVpi3z
TUzUnp8Ssb+ucsVwbQU2JrHQ+ygq48f+wNEK92RQBD2YtnEN71s8nZiP9EbJcHJY
7JQxr0mhY9yfcYZWksEGUkWHhMs2+HM3j32egRvZUrBl+W17SGdGsIMx01qZSF1s
dc6st1WWzN7sUu1rC0F7QBKM/gWQTT1buKN6qjZUbZk1Mr73bbTZonZP+eQkrTtH
4JO3V1Frk2IAY7s7VRvKSiRC/HcI4swbIKKTka/lB5PLDtRZWf/wRsKh6WipOMlw
1Qs4ZdwxUiwRw1aTABiPyPha8H+ZkSz7VJsErCBPnVya6gdGqkALUWn9Kbu3PRKZ
ilq3pVT5hajDP2pe9ED/fUrLxSH/JiubLDz07j6prvikoWQwdD7MHR26abm5bdl2
3rtQoOFHtIvapG2y5F3N5Pg7i80G8KZI5uCSNy8jMW8/XcrA8LXnM0vPdYRiAPf4
/AZW74YN7YXek8U3tqtK9GeTv8OmVE5tQmvJIeJhyqw0iElilq/gFXlTsZ5oYbBg
qDovrwYckbJ6xImsZbPATB7jpzk/nQ11crGNFtHWlXDceWWq0h5BELUN1/bPdUSO
6Hd2CMhBV4CriB0BBywhN63lVR7ZWD36BLSoQLvFP6he/IST0UhEd3d2N4g6d0KH
eqO4qc6hcJOcSFIGSkBgEdgKjU2HRzKFVCb6znfzYbYCEw4BZUxKp0KI2xm4XZvZ
tP7Ot+J903InkYBpKbKwx6dbTSLlJC0bXWZTzntj8Ulyd32GVOVU/7AR4JC35U4D
9e1RTgiB5E+Pp83BNy1Ld2+FpSrlXIs8ZkKLDGWHDyZqS82BFqPXHqiJyVA1rqsO
DrbpzrZudpJMd4jchnGneqXqlEQuk0RvuVDEycv9M2CIhi2RZU4GMGjmqTr4eynG
CfKPmAevlu4LJyFkuZ0958X+dpOynFO++JjoZoRKVYy2pUmVr1+T6ygRVb/tzfby
wLtTFZH/2JwURW+xDCi1yiWjse9452ghOgDetOmsZcvJ29dA0qPxXwUN9S1OV6jd
zIqGtmy3giTri8j+G+9PKWtMSzyvbYKvmxo2F3EoCPb7CT2Ey+J2nQEeU4umLnar
KzCETAOEYdSSlhdjAuDxnYeCGOE5KNlq4IBs5iYOHw/ETE0AT6LHNwn2PCBak74k
34F46FCq7eX3W5G7xOUd+29Q+wkGGDohU5YQ9MxJSwqDLikgqkvbpDqWZXSy292n
SnFhBhUaQpanJ9fUW9YTWrDZ7ZSSVgoM2YXU0cZbwk1R1RJu9qeKMX+J3vEaW+c2
iSmj51LGNqZqL+KZb4WUk/Jq7TBmWL1mbkuMwFMbMEcpWdTzH1YVhtlcWNHc/waf
TcEZUvvuzstr7jpgXpoMqVaj1fbvlVTb2Wgc4laXR0aaPk2Mg0fWkHleOZkb0ysH
1fzuXd0YEuEfDlD2MkSFMG/bkOWQxrs2jYTx0AFkLSmRSSMR09w5hrQoS0qknw+e
Hegnhk4CnszttG00AC8BRPFX64EBP65QyNU7BEUeHbWUWlO8p9w9kO/Xx9LbX5IV
UrcBdWuDGCkcW73mHhDFug9fRHQF8gxRuxgYbZWsAxT4AEhS1A9mgEMBYd1zC48q
FYG1TX8xyS9j5keF69JvN+nHZs6VbWfWZJFfaqxGbejcEndo240Kn1dGRyhwf6Lv
vBa3D9S33jnFcWi0PyEBdMmX2D9aLEzlWTsTelKVtaWl799zVss69V5amlm0gXG+
h5bcWE5ZCcs6ZWWqvEG2xCQXjXfiZri7ow66sPoF4gGCRBT/01QQbafKZkgD2GrO
eIaAjIsCxi6QolJspSYG72coZDawaawrbdv96TIdn/jTF9biOEAFw/TCnXqJk8Rl
Br55QVhZsw1aJgvtH4WTlAzx7YyP3lfR7RsP19+kDLvvpLX69HhLcTLLTZF5iPTS
Tchg7CvlzCwHyOn6BjaLToaZscdpqqmrfTD4rmsCR3bUGT5BNxDoWQpRLePwZMlg
dbFGgLN72/xUhUd6GN/34QOV1fyiPI5b8MpasgNAb6fyEGjlIW3x7q6YOl37eCBA
TQDIuo4iHL+rZZIbonob0jivRM/Ma9ijJofYELOG0kY5tLy8ywBOczXGwYMvQYll
8E1Oxl8Hn5GtJnVyfas9Q+0FDIeyKbSnRibiOztAnIyGp4BekYqIt0QPo9Gqdoqj
7nMyybm6PSpTwES65Q1zVpiA1FfPbcXY/ASqu6Kw2Vpeaab1GwV/QBeiKAz5t3k+
ypjfQ7kx9JA0Jp4X4sHocbkvssaFBBUh296pLNWq5mvliN25tBAmeSReRplxg9e6
Q64tTT+KqakTUfdgd6TWTjt7DuP/V76R2xPEBkCEffiIqmFid8ftN8b2inYI9xbm
oGimqcTsgs+ulaNb7Z5dv9ckAcyaEYCBA8qS0bcXDrF6hRNK+xBw1XYZ+OvjB7bU
4LaIm/7J7VgsaZSDd/cOHdUrPwvypjklBBv7Jl3FdAAVuP898M3OJy8MCxDIf6UW
yLWbjW3hsKFXsxiEegkIZFbaTmxP2pUElMQnpV3R/OYAvbh2yowI1i2rr+pCOzQQ
Q/W0EGb8qVRsM9Os7/Uwqwp6e9sV0qM0A5507Q8nou5YXXKCjqbo0OaKI24wgmyu
RI3cxIiVDfWn8JZKR7/wFgumTW/I3FJqEAA/nl80C7LrBrcKqttP1V1hPr9tCzy3
yaRb5DrGyN0Z/0TjaprS9h1mQkQP+lkwrfZi2yprjRBHCoJL/+3/JosRtmNPOQou
Qw+Sl1SaDHfLpmHMLNjvooyNGI1CIinQWlnkPILrP8zhlMfcmtUis9X7NhYDVQYT
EZFh8zKjLLWcxJGLrw5AhilV0DtpB1XLlwKSUOBSxmfuOqwBQY+LntRMQptHr5JF
7bvjYHm6jdohaHnG0MIYmi73xe17TCC3OrB9YTMzch3K93tPuQgaGC8uyWtO9R6q
7gS8fKdrxJMq417jSqwo9BekH2utPsBEzX08AvwEVwKron7Wi77yGZ8s+tO6SN1j
yL3eTLDJnXiu/3PrEKQOW0NHIeYBy24Yg5PCro/I1f6GaTHXHBbdwbVcUYgYZ+2W
qbcGDlWEunaBIqLvGc99ZdsueXIlZP60sBgiiO2yk6YX/wQGHpxKA2ZnU4u8hZWE
xQ8zQN/BVcekM42mbAvGKZYynaAxWiligYRTalZUre/HSGK4C6lGKPUCTawT7xl1
FjGMimwhpNbehrrVVE8eTQbiz2CVSGpo/QLBEtc1CDRhPa5q9FSwBm3Gkbz9JVTv
4LBqPQJd9A6uErG0uSg7FHlx/khS2hweLSBIOBfZXT5w4BWZC6swpjweejZkYHXN
otquR9HNMMVgpQqS5vrmjU0TlbV7FkKgPzsA9CK8kImJPHb6UPILRy4R6WeRUJ8M
5pWLrf/iDn7hIywzxFwBsXToS/Gbsf6+8WALcgjbPnBkxeZZ2WE9/lDIga+y7JRm
7BmB361s/u02nSV9+881P5vFIyViJcyKO6ROqUVOfpx5W7kdXHwT6EQjfSjfS7co
2qZWdJCwrotq3HCMa3D8sVGQ1hfCn8bZvWrSzwcK/swhsGzZ33FNOEpKu/2mgVnv
3V3CR79V9mkm4jlfmEHIFeJBhffUpbx6gk2lPVO2FHs/H2obz2ua+tqB0+vf35rI
PnkAUMa8qfKy+8cZ3DAyZWIatRlpmWqqHAN8K7MZV+A8W85qjlTuqyJ07pzH5kUI
uwxi9G5okKi1LGx+UGUccYFiOcRMqxW04mmPEo5/lc8RtvIps/a8inAiaXQo2PTh
3pKWkNr6RDFZFhZ7otEEA1cZhGAn6YkdL4RlWjyIlaaer3GB+x76Bz59nMGTH1WF
9uMEf1gEpywj2ixEaNigUSa3aSJnpyH97k6E63x/a6yiakCCUtss0XMIhiGTfwlC
sV3C/TOilLXcK8m0y1HocWINDPf6AiQuSQzcHdlVNQSOewJSGTL3ANVvXf3U1Sr8
GeoIRLYaTxpqx4eYTUAnH6j7K++l023bU1XFOEq75Cyl6/+LYdkyYO9z93g2J/XH
KM6BxVrPbrK/ze38VXGQwLjo4zxy+rRZCUhDxPfjQXlqDq3V4sdpil/Qg0+EW1/5
bEdNFSlmVvrflGeK119gGKBufLgZ9XOkZHCekosbhAl/jMu+tzjRcesTVB2hVJUp
JfzSsEPhYS1CpL9DlJEK6jcRvp67ARtKmfqFl3ysbo5uzMus/QIKroaDR2XUfUMN
RzsOGA3iEwGG/b7CNLcAkHCgjimCI0tX2miw1K3qNO17/3murp+7T+HPJUM1VJkG
OBEmBoAgzZZWpvmgvQSWYrXQp4GQfcZ9SDzXO7kvu3Dh6dEt9B7/RnhHAw0Mr97s
qlrBMIPzXIm0+UirYcm7nfoFDdkJrNXbyHRk8c3WpkaXP2oEj15XvRzF/TgH/xyE
B/kBpBgR6mVppU3Wv3m5uGQFoanD2SCs/VsdXOhF2NMKqvxO38tkKWdx/lkXUuwq
o/5cir84BMFNnF3GeMizczhVMVGmLsIqW1FlAnO7n6yToMnG6C+ydtmTmRw0mF66
PBMUZq5uWso7AIlNbiunRspv+mcwKs7cnfmnpr4DiqlPM51E1rzdXIzhK1phAPcz
RV5hoQKaBf4UF85Wzmro1nBMCKIaqNXAa2aXbReThLcGMTxO0E3drCK5NIgE1gsY
f1ZeX8AY1ONww3Mb7kuzIDNUOOiqAUJrSQIO3e3KwgC4ble5YJLCLplftkiIc7GI
5Q32jQu/vs7EA/rHZwW7BrFco76GLNcomi4iUodkdgknRU67KAPliFykcvJ/WFTo
dKfj03jyajSVeHLgUqho7c7Gu49tecqc+GnNz1o6Lcz/QkfSeKz5a6cUIsOO88+K
jXM5hWj7opoZmuplfaPOuafOkCRbJTH6UyLUVK/AEZwehtbEXfFx0umln8vQgGO9
qVQq1+IdM7c3h9YIVVb4PTWT+g3GTYya0CfYQ2Kx1pV9uevmdQ7KunkVLZZVw+La
hSYIwgB2SCigvg7w+Mw6OpcHkZhjHWoeG8OOgcSQVSbfiM9uAbwOv5paYGGKWUmw
3yDJQLi49ObwBh8o/yIAkW5AdbhPcQoiDlO044TenA4L3MmhsseEk+Hewm0shp8Q
Sa+2I7YGvQ7yjbP0IfutybIK2SiC0SojjzRq05awC3isQgiC1h57Vy9/iyBG2/Y/
Yep/0g+n61Db5LeKQGTqAwKBD5l//N3XcOgGoV/xqIxe+PnCYSsYFcpVnWoXHOVS
OO9YzjkkHlLfzJVW2Ra2TQe6hMu1i6s/M3+N5PG0EhGNPm1Tz/ZvRXFjsIasXpZB
qfk9zyPXu0Lf3Qpa43r0MVkN4lRnv8tr+OoAJF+vfslL3H46FN4l5KPIkqFHarBH
cPS1UM9T2N4iUfJrPppaVZhco934YLfUYHTGRE+9jLvyuUUCTDWaMHdxRDDVrdfR
C8g4wDmdJ03qUdQti2fcIKU9Dt4XjGB3aawiOQlItG0aS9haRIlBn0ggXC0/tAFo
lvO2bokia5jVBlrFAhb074hOp3e+hTxtHHJFDWPIevJzUx/NKxkjRCW5T6ror9nG
WcrVjrT1Ffvfo5Xwt1wAIlt77nR/HOp7XN54SRbEdRJEof6xFLgMMvUN2fVnuV1D
jvpi0ESb+YVaZstPOET3d29ptjCI5mQApBe98mRM4igxlXiyTnjhZQgkLzIilqgT
xeMzCFOJOK7r0uEHnV6CTd85gC8jtQRLYpIuoQziwYzP0KFszB9iyWlIqBcmaG32
EmJsFKL+Whnd5SUNjPexpQO4TAuEv7GNyHdgXzVaSLUPOOgD78SiIevF984C8uLe
ASu6TxHABs1Bg96Hv8DSF3NpOsIpfpkotH9qtFKYA2tbqMaG5Yu15L5xu+DvTWcQ
49A2ZoKyVZulf+Iepym1slhJByOkAXbxGYx2yo4C0t3QNVdjf89d7rf6A6YVqDcz
3zzkTXG3/GAEPW5MCwB9wjPLKJKqrVBC1+ZGB8fj94o=
`protect end_protected
