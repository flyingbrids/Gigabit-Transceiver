`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
SewlKs0AhtAx+77sQN3DNKyT2kD/JAJOt8V9/ykEm/ASjoEbCI+BagRYGEYKwp/d
alFKlajeXBiiaWE4XbCM8VVQ9jSjt/o06oVTxGc4nSQEz704unO54Ve6E/GMsmHh
HosoR/PzucFEIuVO0RtN8Fy0Tku1CZFhqXgVVNP0BMPa7kQLKi8fCnFO3tjthGCl
EacIuXS0Qpoq0cAHsqTQb35Lpiy+fYUuiy++aUZ0iozhzLq49rfdp4etL/qt45qR
zeYfmgCAS0wJbHPjquKHwARcc0oHGSEqa61vULeS04qZwC5rAjOxmGuRHB47KC+S
of4zG3aNPqeXrwx5YxTpqA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
L/HV5MVj9+DtNXqKJtefnr4bGWviRmuCFRSWloJ61yH94FRgCwZcM0Q57JK0gzgR
iLbeDVDAkQGAuW8C7wsT+L6rSi6LQlRpJCjFIV+CzOa6a1VTE3WOoVY49a9cxJuV
G4hJgeqjHOmnIR+uEWyLUwDQw8sBr0PPfMQJjf5w/YE=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 90704 )
`protect data_block
ETD0+PQ5YCqYl6BJijQJh4L2mu9wdk4kb+AaKwbGWVFxCFh5ZwKxXyyptvlFz5jq
PNHomzU5ZWuyow8tMvOefM0btO06+W4j9igMi5Vw+Kd5EsmOnERsSVTduXU3v3e/
Kbt+f3oZN40nCwZf8gY2BizQSixrFlmNyInsCPn634y48hYi3/e9+tA5xD5rUeot
RWCBPWxH1rhEk9yh8PJ/rbc71g9h2sPWNxZIYG8vtvA0gbgJo70AUpNztzZX3qi+
9t/x0eD0D9OadpLBHGGvm1X6bTbR4fdIUeQl/bknRzbDemRYxeFlHC+9O1oKf5Px
caQc6dINTDIT5Vx4Vsg28aAi8eS/EbR2YPZnvtodph4lNA7HN/0fLEf3z48kXhiJ
o9Lpy6yR++xBBimZpf47VgL+KpwX1f4m1Q0xatcL36X1CP9K4QANbyItBOi1k6i4
ZPW1pCnIpCVGJxi343t/mk9Sv+0hy6v94lS3bpNJSJC534/SGyZ3uV8F73TSdeTH
ZJAiJ1w9SPbkUBCbZL1OoV7Ww7/0DLQtFATGFuzNUVaGEMiliy6XXN1olH0bN8fe
T6UR5B4Cwv2y3OVAttB5pEuQbakZ9Kb87okbjAa58LIvkcGgBAU6PIkd9fq2I8Eg
yphiFaADXMsmbIAkG/n+VlcXUAZq8newmERUmyUOxDbFQZyqdxbmm0AxWAp1qOD8
ZPB2e8AP4fxAc686ojkQjYKB/mzWGOYXUyjkKT84Qn1OYUYpowa7susdejfvQTHU
vb/jTbtaCLBMaDe4neLtyLv79PNzrhH0DbkZJAfCARPZu67ORoRaJfpKgJye1PkO
J5sUmCv4byaczwj3IwZNcpmhuSHbFXJwy90dVS+sPN55J5f/nmRwRhyecW6vMWSX
J46fs0fynr5qB+C2kg+MHicepHIUV56uaH4apyNQiQGnmzOzVmmyv+gC7oM4SZ9p
ZcKQ98SwUHpjMMoAMgVQFqIKrtGAyAbl5zF7flNgZ0D3ZPAnqG0bss7a/uB2QqTe
+4bDruOWwh/iG+ddYKn2LVxW7UPZyNvSn/PEMXZ6pjqevubdJEG28qIgF2FFeDw6
6GxyuWCdbqzFJtwmN1FXeOwxmvwsfZehBYWxIVTFTKO4iLTezCBErwpqeWKTjiyz
UKsIAXeWlc5T+PcLzCkyd6ARZds4JtzHmtThdrQWIhszsSoaHpALp87AdQnt+bzv
1ckixzvDrOQEDLLDmK55B6spAuQ8nwewiyNfNDjoNf0/HspkkyVb5T2rbzvD1zoj
BfEN6052r+7S1VtCR1NrGUUf0j5pR5jmWDxCmamgAl3OPESbTIhBrrPf5kIbJaSd
Y7eTyIDSdMmZf5gLxQf+PvG1KWP027AwqMNWe5q1FjiEaSPthumeXbVEs+KdrE/r
rqzUvhcwSxg1odQw5BavOE2ersvH4y4ycTrHpbOuaBAiDk/LNQaHZCxsQnS5b6HD
HyFH3Pwnf5UVDbXTQap5almr+PB1zoLphdBSNPm7wj7ar7dcck8XKFmvooNc6DL7
v5oguew1prkJN3EH4qtgtCbDl+bkdOAgzzDUUiJBGg2cBk1s0fMeyZnLWc4h6CCq
XcVVrPIVrxzOlrqP8Iv9aiLZgsInwrGq/4V6XFgyWLFwbHuKz9pqJqx71leMXCOs
oXKJzte1EaP8OKf9cS3heATLZYFXnXYZmWUEjHS+fKkpgr0LWogPObvWOogzDsMs
Zg7jNCElKBERWys+Q3dLDUijpRspMMBVMnFxFhWoYTcu9gXDRHUhmO+dnYDjJaUf
NReqOoTpIuDvt/grRIn0mg+ul1chK0ebuGLzRsgsav3cMqgtPMQepRrYgnNBaBaW
CpASUvnYHqPBIASfPh+WNOBaGLuNgWGfvSYwRVwZqZErCKThinYfZeWyVfz3ypYP
Z0WZM8Qr/PAUQX3td/V0FIHbW4Yg2Lhf1/OYSl+zbg9yN7PyVfulluixM9JzcA2M
WnDX3Jc9vqzH0nkOZnZcAOlh8ad8H5KfJNsvEKPHFSd4FFP5cJ8Y/pP3n7pQ34DR
0dX5ANcAfy1OI5Wgvgy2kDhzwEdtfLc9Jomou0rXg4UFOPcDy+d+cbPfTXcEG/o/
2Zv6/FosMG1FyBPy4RLngKhY/wZmzBRMUWldEpSMuNbTF62/CReXfwWe2PnyMQd7
+rYLb6Y/nbraNMRI6WoHJi7BoL7F9C+m1pEK5AMLm6EAKml3JZY4jkvDt9F45LHx
aPH7mdhU5fmSnxUcGGUqRQiRP62G1QR9Wg7VPjQMbc6l5BLnyIy61JeST7dtxYGr
sYd+eb6NDG9Gf1tE9jzM5GxnIFvUJi5Al1UCuoygQTwPy6ego18Y6VA4AnmiBVbL
pscF+X2tEYHWggUt16i7Ff8HGbxlIrXM3+PBrxeU1UsonWQoxQ4jN0b4Z+YLcyXI
OgVDFGLseZT0WaEbGTh1ezscz8R8PcNS58O3mDG7y0tTkco/AejW+BLlm2NfUMzI
WSWwpZ1glJBoXYzzrt57PRG6qHR5LKL+A9SAiRsY1MM10f/y1z/S2r1ZPQmljOvV
bl5yNjloeqZhgPYPEQn7tR8zOCo15tGw2eSoeCUM3jMbZvN1nMIL61XfyismXOqu
/HNquAh/OApS4Lf+tjhfasln8Q8JR3IDYkCMRkM87mrCNpe3fSGXWYZ4Qo8i+kZB
mbAtzLFu0u7wPD6A6n1YsZJQuh7rYbYiEJgtGEm0hqskigIgM36zgfBaarsepcCf
b2zVjeyILxr1PlN+5q+WZkYJ4ryhLur1z26YL+dd55ABVolm79csGU0L0Y0qMkUb
CEewla/un6q7ODsVuYhk2pV7u13qiqBFIgOCZGUEeVBwpEDAHbEaXDh77M2A8taW
N0RiGkKlwe6oOIv8jRYDM5W5w1CBYysgiHVJI/i+bQ8ugKN71CWEgiwdPVoi2Iow
Isnzkue0r0hRoApmxmRKQJzC9m5ZA41blTXEOmdkjvBMFHji1v3z7ryq+3+SIdw2
pWNQ0uYYP45NYHLCPAMkWA7xOHLjO/0684Xw04Flx+6+YCiF9kXlfT3eMB6b08wc
H3Ey+TN96r2M2Nuh3y9xIxsWWoa7XqoXo5VHvrVMVqGRLi7972wztDUWcFYFocSB
6nWisjK4MOxnIOshXJ8fDcT9her9xf+0G/hlqYTzfvpQb8I5dE5UwxbuA/+Tr1JA
P+HXkSMbFRwRgsGyKe+2wpk7P8FNTItMhLy3xO3vEivCijUgMztqagJVs+ujJ+f3
4h0pCAhAXzK5qYyH8Sa5zhaodmaRKxlz977IsMpy7r/A7BlL9VJfkXhLJE7onfAy
CaVkizKqgzclBuqGc5ofzp0bK/sQZPKg3RlOWRjlkV8BQhnGSnRKhcSD2Dr0ZiR7
e4OvH1IgRzkU/BhgmCJMDKuo/VdBSpBDd2VjnDdZUrqRT4tmRd6jxdYgCliZRXCo
FqYoGfRn6wGVIUnxehVz4/De54C9BxhBOpfxkq0wgjRx5pcRQDzJbEdy4clYJLQK
Pu8V3de1uJYsED2c+GC7PUm2lxC/GyriGgoMkezV+R7vfUAJ874n2DX4NVQnycK5
9el+6vc0ghZM+dXzG21PaeHFwRrtraenHwU5iTHTQEMGZxyp+fLkfK+Oz0PrZFQP
BdzOeTA6xSAnlHL7Xr/ebY1qwhnImlo6/U742prldYnFvV9hnFAj+KA800vyGcM9
VQZ9uBGlWGo38hMRYJRfhUKAzMJPe0Anp2zWeVo6Yc3jgftLEI2+Um96mvPGgkAe
6twVPfa+PoXux7paTPEOaqU9gUEEFRTi9AheQ512aD5yueMyNcrFvww/NMqG5m5P
E9x9zSool07S0FMLFdFOSZbaBwag4q6uO+e6rcxIOJWJ5OB+NJbN02PbTa7uXJvL
xrBr4wD7X+C3jpTwuqW6SFgq9uE3SOeTKxPS/LUsBBBOUWA/lrXG2pifMQL9KbY0
AdFY6T+KnfRl5E88ElvCjBrF6GWNJucR6Seub/tgKrRfKGtvrJMBRMA+xPiMMLPW
h7zDJKlzi+TvR8RTGnt3r3Y/JzPloAHUiI+A71RZyphnJmym9al1VfMP4Q6Uy8WK
cP4KgF0S2ZWETmuWfKPzH5mgVttWJEF0aG6b+xGgmd925P9E4CTTyNELk7H1FML1
++S6TUeANrpqsMb+fBevOv+spPHLzNqKYyZ8dey3udvE4LO9VIZmya7nGj+zfHDR
BawYVhP9aw//+FbcwgHS7Pq5GPYsT/le/eUvDpbyOfUCv97MR42pChslcVER6pza
8kMu8YiY7FQKxxBNT1kqays8XNwz4sxwHqBKxBDYDzT2rHLA7OXowXQgE8W+0+35
jHINadiq7yfy/gn/6Rq5KSvbIjkzBzaduj28sPK+WY5M95jgXj5hk+au/7AjzGU1
X+PGenszzCwC7+3JW50z75msq00bFzd0/lpUunrNOroBwAxpN5GAuDk6BBp5looJ
0lR/cGHl7Ky89s6jlC6leIpgwXS4UQJVqTue/uzcY+wR5H21Ygt+5rY+I74j7o9k
eEOvX/7YLW6nE0zMgHRZ5Poid6D+aKG2yDnztSkEWXOAiKmRMFa7CkeMVJCNlAq/
g40iuB1IrWbgh1DRPEP9ER9qkAhc70uJr1TctQ+gLPDegbmBuR2rB3y5YbE0NFZY
UpTaBv3c6AQgWFixEqPEgzhUX3cYlFh9kMB4HAURBy2NchSpQXNBqIx4Kp6bPg5Q
D6h6Y/Yf25tU1TdvZJELL0RnJ79f9ZrKFDydOrDGxV8tF7eGKiYf10bBDhPPZtpz
zme6sgd7XVd90Ho+5tr5ez5hBU75a22VM3RJnbFJdVgHjP1J6iLO8yrsFQ4cvvxj
Fi5j9702HsaNm9fuCVK6mepi2LRgFInfWZ1fPxc0+cCEPE3HZwCfksx6J7DVsGxY
7mZqHzU+u7GfM07LbI0xtzPSFsFII2ZPhMKedFV/8bCmxeCX6pCGjQMGelw9sx+8
FawrkTMtzIwXj9CyPdAGiwJQ2zwEsQHbnFI9TEb4U2dDxEKMuzh3bPLahahfeKLh
4WuV+8yEbMD6pdumWobArzOXTkFUWmrM281mlJKV8gnWRvDpHIa65ro9Y8r/LJn8
fE6yd932P4rTMO+v9657glgmTRhJIeIVoGh8ItOQM2caHGy3/3iszR8v3nFdMiby
sMIMTS7rqEyudG5lX575EsjfRm42UJpx9cnu0jRusaJja9qr7fa/fjuho52R0JHa
1F3+ZDoM/wsKwvF/7xyn5cKfPhXQk3oWk5Yx/HHi50UPuUb8VDAVar2/UKMm+yHC
jjn8qKZLRGGs9DpyOZa0Ak6KcxtEPWCjrHbF1ICnVSaxtNzpUHTaJRWQ3Aimgfx8
phxLvynDe6qPsr+xjnRK3EyS8QkEgR6CqHEqzd4gEeHVoMb/E4rCTUUZa9Zto3i1
WJoPJSZkclKbl4PqqF2Sgo1EoQ7yIXlduJMO6RVla9DdpY5WdYW3+04A2KGqfQyf
KvW8CczF97EGxwDWhqO+85Md6kECKu9JhmJ99qsF7EHtD3irJgvXuswn4/U0Rtcp
nH8fklZppnGx0uJ7tCP8kUYuIAS65uPZuG1ZJOD4xmgHFlOG2zZe99rf0OeZ934v
47t5lHPXzWVcJFtR99LiD4iZbF2/rYFZb82cyigjgni+4ABVXpnYCYmiPEWTMq3I
S4Zx6vWFo7pyVV2NPOWDy5PQ26rC6vcR+84nAx6ANpjSBXdVtI97NUDwkFXJDd1G
8tVQ5OeEGtUJmXqrV9IdJOARHanF8FKb7imACCz4UX2Wc+0QBkKOIKGMbYvghGMI
f59dz0uMiIT+o1ZjhLOqPwzz1MaTN1yS8ZKBc2Kk4JfN2a84SAcC1kDtYvr2ytwi
ekBW+h9aaaX/LGntMmI/DrnCzM4yL+nt+deyCiNNMBYL8up7FB97g4Evz8imErki
ztTpxlMJ/eVS1mZDIAkkufG+1ikFHYhYk4igRNzNY7tyZUuXnGySTJlbuRR8NkcX
2rsC5sMAYq9lRCzk9B5n9Rm9+/BYHiDhKOa6sSt/Yelph2+risQdF045rexOvoY3
0jGrBRj2u1DPqzvzlUJFoSV/6cF+EvTPGzI1QnuigVbxwjcwhe9G+oFgZT3Ku9XZ
p30ITqsXcsChwTdp/csykbeadZ3XYq08Xq7QqforQV3dMiKDbzNVewBpTz2alrnA
4WFvnQqAd26eQ8XQRhlNrEkM4rYpATTk3+ixtBZ9zwg15tGUppCTaXs/VSside8H
HngeAOqsegDK2iZD1LfhNEFqhMCc7Fe9rY5ZDMGHDjRbL12y7n4SvVcSTQwD1pcI
2Von+91HQ190jwk7EyCZhky8VaySgH0HGwLUQYI8JlvhEchbFK+Warm0BdCjQ+PC
EIVo9OrrvFKduSFc5TDdkKdqFEZybnufeIebP/oqvXzx0TS9QRUEkPEAq+WExrn0
Gd3fIWtpgsyCVxvbHeA/WcR51dYJSFNrGKXbFP81kJtz5f4XOOs/8RweeFdjkhDA
E8KOXLvbcrICdKjcqE4fUHhwTFJuEv1NNqLNvkqH9m/2H3038hqdR4ro3yeK89Uc
ZRPHQG3FfmYTs5yUGz1+pjDmTuuqtpkrwM+4LnPusu8y2V63BgNsq0mWk/CPao4/
WfeioCor1ZcUFqqiGqzV7tqB5sf2j9GB9wxc/GwaS5TCYfQGwSTx4fb7y1CI7Hb7
Ajc3PC4J+xSaBf0yvL36gDWT5KTbLPCBgZKGVGf4oKblQ4Qj/CopVlWD+QH1oSHM
gfh/Y5efnu8ZqHXQjNATnzw0e+PWbUxpe7GGBH/QZFFwaPfVHYp9Ff6LljHbMhER
stFwxuxbSM63rNM3EhhrXL4YAsB/jso72FxT9cSLAZ3mEzUpUnn8BjXbO1Gi1pxd
0+K5sBCUm5h6kCFlZofiS6kBHk4JQGwX9DhtwwimhJhq/Ugcy/s2/F1u8SG093JN
eAC/OsDjcZvdXRD4786VPX0Vwty9mdEaZ6RIW1LLY2QeLdZ+RElWZUUo6ub15uRM
KTxEpYMayjV/WDaJv/TCpEJFenKMYPOg5RF9INlj4fkTKy39iKN8wKoJNQH0GIDN
uaSaYPcgj+/2yc1YDYsmWE37nDJL9X5BledDELKShx4iKPndkUW0wH/2gVvLUzZl
f9dlz3Nw+bcfqAD5aR1JzlWMNqgmFWr01tZ4AYsphSnqyJpLHe9SL/eCfcKy1DR6
eG3UwhUVNY49vv4cJ0BXBAaHuK8nfUZt+iik/0etgn0/IVKR1cwvsYh/uh+H4VJW
eBxtTfDg/9XfUhr7q5DLXycC5PqsUVBc4O65Pj9En1J14pSJUeY3Nk6fLPHCkHX/
mvXe1F9M8k/UKqSW3eI/LWWKLO0BmChs3pFt2BMaA9q8YFjtk7kohj3eMlLfZSEj
2UrqdCLzFeAZKoK0hfnqOSlOP3yTgH7SopyHjYCpJ66hPr5bcbvaI6R1kVtynmLZ
dH7zWzTq9DHEqvjil93x5pFdtCDxrXRe2Pssur5TuYkWTUUbWNbR7ZLXZzr4MvJF
th73vSCuv1ws4OCTA/Lncs9G1iGWIX8sZ0WTESbdGFt2qztWi3VqXhd2R9GKQzY/
jtUBJbnQcOa4Ff0sRjn8lsJ5e8uMvfleT56Ta6JdlBsy+J/Vn6X7IhQi/OOUyNvR
cMJdvklfPAVgtLbjU5STIwIZ3+OvpRM+4Ev+13M+7SwlcDhEeJU0BJTkrP93iOth
qBIiTNnzRDfaVYEXGVXwj2w2tquIRjv5sdpNSMTnStGanp/W+m6mGMdcstA826dg
0Igzo93beeseOOS8XjkK2pKgeTI3FWeC1jjWbm0tcD7qth31ChjtPZzodFSa9xCT
jXco2FNx4FV13c/MmM3LcbzPvbOxoMRELbKO4Agh8FkNtbQjEYOeKJ5eFifr1TFr
dVhWu3DFJtXOD3GYqcV7L7W+lWHM3uFBbHb2kfL8c+9jQdfJ4JwQjuY9gIloJNwR
2ye2vTVb1W33XHJkRZDAis8D0Hn0tpl+pRtLKRbkdSzSee2oj5dZ3eMioZ1ICSxv
eQKShHeN9F7ZY0KQfd72WgQEtqFr3eAHtWH/n/kuJvALD6GQpvHuor5j/Tph+qvj
n7kXQzV9jP04c10ixZcrUFig6B0p0w8RP/VDnpM8jZgCsIU9o9jjMDr39kTwFlFh
N4KYrwqJhytT+9rpSwY6bVQoarq0OTwLTO4rElg5KsjiSy3WjsKAW+I5nSMdf8lL
qT5SA+A2utodW52gfoc9ofVTvrIbkJPoOl9wx++EBX2Jjs6UrVV0o8bY8/cIv3uy
urDYsn6RF92b/GlvsWUSumeCqhJ95LqynfBeuBGuszbXxvkti87CF+XbLKMxIjP6
Tkq/ff4KXNcsrFOB9nEof06YdC91EGt/qtw8/NGQvV1XNCAIEjckp/qCKrDHKAAR
6p0hG4tVYqPVpZ2pspM1Dzi9YKN/aSQRsf0JiBv/MM/rnBE/S23grda0l0ty5Fa6
ubOtORloczcBownkCWzB1+vgbeYlS8RPePNzvQfONEShVtSa1L9Aa6Ji6N07VhT2
kmHDei7zzdu1VyVnTpQDtVeDG9uaIbzJtCORUTdrrZ7LRzhr0+NRZaNPLqKfxLja
y3n/e6ckzRo6LNfWt+ufuYv0F8GEFJzq0kXT7BKes/8/NkoR2ssmZIsswDcpHt/S
Whxq22rmMb7/JH77xB7TO9m+dy+0jjpPDrSQeH6Co/KPo6Bgk74s9YeJ+DgI3hRk
zBG2mXqIP3YD8GkkCDotgLHRdhVfEMmx7BiaYXc+pmi0r53UkcfY00TQ4FJSETag
zmgzZU7c6q47upn4HLqF1DEaBdndlgiSgj8+xVg9e8lSdrbSqiqmRWrbUQsg30Ou
35qzP7iF1doqad7XV2CVoNr65EotAJEFZjewSsg/ZVsle6JE1EUAamvtGpCoxuey
hRLF2RIf6IGvEJCtSuPMFJJ81OKhA7X6Y12jZTLQHtGD1DvYVTNo+CZ1YC9kr+T/
6l6NcofNemWJJpRfmHOhWzS6TC3pyzwUZhyp24SPaqdHun2UNVLLdvmFdhFBswKa
XKQXZndIPbCvCKfJv0lYr/5RxhPw4wnQTSbv3wCPBGjBiAwG90VMXRe6ExLL4wno
bP5+uhauahlcNvF3mIZwhL10wIQngVfwRRI+05xl/IRrvb6Xkej4VucqOhF/HsAN
zz/ykdq7aaJenIIyWtygTADCIkzxXKVzcz69LHRCQLyE+5EFB8HqMkAfP3MmTEvz
fDhGmsQTisg4gRvt1z8V3SO/ZaomLULAzxaN0V55mIckekO5lcBHRv4SEoVmDDZo
Ty2T7LQt6rFioQ3Bi2czwnfV6JSKPapKNp85fwEx4/d2DM9k3Ey9litLKvh0LHjT
OUKxNRJQnRIvZxKa7YStaXZ3WKKGRdvnrFXbul8XZ5ehxPLpDsnFuDfRTeO54vgK
x02lscSMk3heIF5UEqT3eI1baVbXDvXaqedelq1UThrmcMhaJLBrX5hkzeFSfqVC
AoWo+WoGPO2rAjIkksN60pKcTz6+YLw+l3sMkUL82ZXpLU7HY7sf+thqzguLCaGy
iKXZcuAX0OAGzTk1zzxSIHy1NUZZImQMRzOoT3qeF3MuIANPxN2g1yx4+WmIqzgJ
p8I2sracUW9DiqkrSqBGe1B42MP+8iqEgbp3IazpmWDgc3xOQj98Zy0Cpm2Jsat1
jUrGPk8xuhQ7XWmrRvFdK9/LsacU7V44Yu3lyJepi9oIVDjCrbU/9FK24etQBnNU
Unu96puHSUZdAoSYxovLwQW7TyRpQNcUF4kg493g/tJCbsXhPWKNKsvmX7BI9Vvo
ob7O0FJgcC+NNhoX6LU2s0/jyCak6XRHdWznlWpZIUouEmEOO4suvOPnAjdniwTS
uZz/ULlf2S1qhlMXvSN0B+GwtAs8WwkbqNPkAK+iY3zk8w6VFM0/6AR8aRBawZHd
5qEmo2Nz8Y4jaJ0fnm4s+a5YudOneYTmVs6++o5eitS9F8ZTBLj2ooPKQKHAAUDJ
3UFBZCS7APnBu0wnQflAb/k2zJPGHQqheOzIYTQFWz01OYo/tCPWxMFha5LvC9sm
YKXjRNZa815q+JYU2trKiv1b+xmi5OBuMiudzRFmYrlw3QLrN5eDXk2O3vNEArtr
tLkVNP+vcYiIst91L2p65ub5qFdEut4h2qOTr/jVQlmcGv7luMjteP4QmtHM4Lq3
TZiLCoEzKiX/ewA/ES4pVKE/QZzK6VZyM9bq1L8HHnom7QS1s+CNIERlfQXdxLFv
F1LrffDVn0oN9Dyrv8MZZ9MzZrdtiPERDMaeeYa8PZs43TT6Eb1QWfpHduqPp9Z6
wsruXyRyPiZ4XiWpF2qmsemFe86QvKa1B961DcnIDpFWzIif+e8SVfD3PutmhDmM
nyBEgkjJ8RSMXYTQeRz+38bG9FR0X1uaQ5oBzRE5V3MDKp/ai+JLy1qsLRrCLHaH
e4Mb6FfDj/L/h6bhffoHqAvKiWjfFe7F1TAcEoTP2tGNhwGmUlz5ucmMT1fsMnPT
n85oQwPDGEe4/jIwPk4V/hvmwruF/XK7ViwfJGglb7Hs8Bd+5BHindv7h9yjW2tS
F3HEh5pp4qr0aQMkeXKtbo5CMRht7unPPZF2aJjoEuxEk9g2iF1N2pmhSMRY2K0t
eOA0UyVCeBtEo5vGFGy173z8xGVz/7ziIwyFOnDhKsNrSO3wdD5Vqwk4YGORep4n
FTcPbU3vSn1cMsEtNiB29bxyVXrUHRb/r/uAbz8vaEvGEwMoXE119ei90w7/Mama
P8GKAYxVgcMMT5+QQ0GbK6FjWaEmWL/EG6zMsdVqkyKASnQnJBzVGA5CI+R/bNP5
1eYQnS9VSoLZEgnfOS86uxDFspErUszANyBdsknGvDtM4FfvqYSHA6ZkMnjCDBCY
/iwmgg/sBC0NW1s3YJSrlqIWRo5ZRzCfTaeY/SSbNnWk0i9Nb8BOKe26YON85T9V
YKvL8Ht+Jhlm/W1NaHk+My/waAnTqvXuoXZ5qJZAoVl4cseHFuAbTdGjvF1xCT8J
fmK0QkLXhk9l6AA9zLa62qCG9BdY0U9IJ9PFzmhxLq+8SK4w8jezsWX86lN/2Dym
FF7lnjU6WKtD84xnKR/9lFHyg7ZfoAqscs/V3qZBRpDWOFuHaOY6L8WrmIpBLn1f
wlp+Mp7ziZ7BuSPEUCzDP2Ea0Hzpnw9xepgJqeHPenUUOvWO9gwGFd66FWfLJU35
LtX86Ej6kueHJu+3e/Q6zwQmvK12r2rOMgxgif3MnkBzBmMUZBt37iZ1LLegSLyf
XUbzi40qN4QItXOwRCV7p/D2zNuCQa242ftbuuOBhkLXjTFvlYMfSE6seO66MWnG
t0830nG2cdyEMcgqt3uQbf+qfGTMQqlTh42Wk/WjuVmy0fCJqfBOCwiTx6zdNLqW
UPnsKqGxunHUAO6O7XA+1/oyQVbI+6kkIFwTtcABxO1qK/dt/0QKJBRpq+XRyY8Q
la9q4NVOeav0Tit1HVmcUj7S+9TPuQg4BymK8whLwoP5MH+80EOVJiTAr5g9zbf9
ETWXrvS01G8uO4JDSB6g1chpFRyf5o5UHFWMkZ85OnDKSEt/fWk3UE3gCMpPhxCv
zXX/n1vqKbM7GSUl6gbL0gxG4EwBopJPQwHWEZX3fLhM9mm81b2KpBJjsThWROVD
N/BbNoX1mQ6ibPARqhwUe6U+yKkfBVrFF0IhIthg4RZKySxFv9mwofLGZE7Zi53d
4ZXvS8/iJvbjDOI93wyxvl115BBMT1R8/w1hjfZbwvj7zvNlyszbxbuUtnOMvidq
ctYPuwgZOFZU7GyY+3MrWLIbKk8Z9McAOw16FYCtgS56Gsq0Oq8H/vw1Tq3bsj3x
VMTVMMGppS+GetbazXIjxr5lK3pGePwgs9aGrQ9EG4BVTa1wdJjwEQlW/wRokTpS
I71CsgePUA+UnujLFZzfr0qN+AQ0lDI3oQcxIKIEgEalTdkWPnQNobNG5jAEUl3Q
Fzk42owyVjCBiK46Q422JMcHcl+l5AHPfyQW8v2dzKyfguzmQuYiiDUJ6yjl/+P/
kGYnEWgM25wJchnXH7uUp4ebOIN5EhplB84+VGFJHPXs0kq5hHSdKEYyp69Vjexz
egeK1ept1aw5H9TnWFO/hUPTFE1ZRWuuXAdP3ZxgzDgNdRD5vqSTldKRHjq3a3Ug
2r3+kFWJysVLa/c73qLph6vyQHfjH9RFWc2jG2qzVpcRB6N0+FsQPZpFj+rdVMbE
V9nAFz8SJTnMR75YMJ5cSPi0Jdv65l7lJnaqrnNTiaT9sS2is4QykEiG9DMVyl3+
QyitrgHvRSZDKR8tnpZ4RlpPts6P3JcMqYtbqkHJyaOiuwoXeFShRYM+4homakVz
7qyxr1P+Zp2hWd5iaKCPZUVITT9U6zSaDrd1/eg3Z5iugFWUljPcY0vWs3Q+18JB
XrrTlaYu/niZPBwhZBPkHx78+YYGbzHzIs7opM4KeXQ8ykbeY3rEwjEzPveCRi46
6wNzSnDjj0TqHCghcCP4SRTeQWH7hh/Uv86scBZ7WgQgXPn0Uj/74cKjUf1uNOOn
vnsK8GsmQXfFcUTuaLm/joqLMw9zcmTcyY4AoPrn0d6Ekl+ppqCM1/1oara3Iz0L
TA/VhhZ5H/CCzw/c73BZftuhWsXewu0eI5xRFa+OQRnf6FV6KMmu6C7CCfwEd5Rb
ldV5HmkJ71MuUVtQDtbsZGzbcNX1BMWMrBXQbCww9U6ebRJfJCB+O/pU97gQi/Sf
2dXBIlShBh2xHmUxaGNPGki7z1NyuwhGH9FhO35Ehvp12rp9AVX6ipMl5VCS2AG1
47kPQ9NfeCIMAwXv8OVcP51HukTGNV1MrPqcCuzMiEX2arAWDY1BAwLAVj3u3dBu
ltlmasvq+HYWdqGigFBOxzXB+6NA9paDUn7dC7raEdYnyO9uuCJKBOjmBoWCFxdz
cSdWKE6PGdO3nzi8KYelm3tyRd4OJAFJTnkJpVVkTnz6so52j32u/QKm9xPFjqIc
KwzF/1Xva9EWOdMsb9SAgdJMwIT50jTmqdG8uZK6eufpOyf1ohNaCoYffy/Dsn/m
NL6FABneOjLHb/dLCZr5EXGjkTlb9foWsOzafe7iEFUj06fzXXX+2sJV0FP/erpC
j02+3rGo1xWoWY4ZDkM7wbTdXoi6F1u2QEMws2iSPDHEZH5df5Fb5zOWTRb8yCvq
I0OaJtJfjERwAlL6oiTg/f2nxwuCB3OJWXoMspu7yTQL1dIl4goEYeS6pHkKR8G+
jA/VhJmCienpzH9jbSB2N8sLBkrXWLoltxZUU1VclsGOBH3OSvI5osM8hs9RK24q
eSgNMuvmQcuWDLLmTdLd/HPkHP9eA1THuxmwRq4zYCQx3uOJT2hK1EQh590ViQNi
Iiay59chOLrPMwUIzmOedvxlp8PnKdHp0Rzr5jZHVTvyeIaWGtMA+ExMLkUCt/Ia
VaMdYEeu26WQCA54SC1sUGMh8F4egu+pnXsjrwElQQM0GrU8U8Nl4IKLT0A3K45k
OHmaYDHuuxMjZDuaETIGOStWl3U/hEd3l1KJbU1Rj8Efea+svlTELQhO2b/tiZ4C
AJB7qaVlkfCLT6lcL8aMHphdGmIGhbmaKk/tu6SoO/JWZe2BZg0vtZoqo8xfLhN2
/i1oiOLOfYR/z/zvdrIIY1QDJjq/9fyznqW06YYjy+93EnXMgiEZnNn6G/6nfVt5
xji9JH33CsmXFPfo8mq8Ja2hntwXH6c2BxYtIqE9iG3SXwVMigC29AqLHbYkGwX4
TUEB1x4mfO71oo6p6bjSj02KOuzGFP7jCjNY5+x5BU20bRcRb/iTnOhqIrMRSsrk
W+Z7zObFvc2jrBifJwqMGjAsKarUCFL26/372ROZb31IePWlhaRp+zVsmza61aV1
WbqPXFSgRixYI32vjjyfVLBAd47zIf4rJwa/Mj/Q31QZ9dklUmRpO1/8ziqudhMZ
f1GzHTBNRsWv9P5y5Es8YDOKAtjl0wFREFQps76y5fGXBBe3wp2mZn+F0Xk1ex/k
K9x+gCGXCJAWFRGl8OTfBHklN+e8QgOB/hQLaVxeODUY1RbGHcTehcBs38LWn8G5
gd7PSQAKwEc2a0BHbUxXqJQJWPaiV7JJhOtmu2AT+OU45203dYa+MJcD/6iP/IOL
lyjmD8QWZepy2f31EsS+Efr42gVy00wJGea1JcGTIml0361UpSXszcHdM7SJ4htB
mwhKawR/5z3eJbrhQ27fNv1vlwq89WCJdkhI4zhWc9yMKluE1WtiPEV2klbBghL7
OlbtKk6C/Odc9BpvCDgJXiJJ5sd/Dg078boWn5hKFcS+zzt3YpQbMfe6DKqGyrEo
XEcupkGDc5iJEzYlI/+lqKTGf6PJLffXW6Fz3P+sdc8wWeaNG5PDiCHjdkZuj8Hh
hOc8DFIhBDhIDBrIiKQQddx8INKm2HtZxQsibPKyxqIIRyZLBuOzbf0mCpWaG1kc
oS1vIXzvwhc+oyE4hCl8YzaRxny0OsFRUchlCdVMg3+/eE/1PDsmBa+kDJEZihCx
RPHUd3eaR25WRfb+d2pS1b8D/wUgoWXEAEEAYQq44QGw3Fta0f4FIhpG9vBEI/Et
JOr+UyMkkPJUKVBWUgo6dIasyZUXssaX65Xu4dtOzly0KiTNH2TJQJrQ8tPGdZPB
7iQMavEpmMeVdVVQ42vVqZE90NJ6APKSYaX7mDiPiB7IkhPw9CPOCv6ESJrS3Zuj
BCQ9Qjo940pz9009IxJkz7SqRZk1rFl0gzzr4DamJnlDfoMKTvhMuZEOLbuPeN0Y
iPZA3E6F7yq03TjEMxPBEABQlKHjlOcixT81p7nLkJycUf0FPXljt6a5sBoOBV2N
v66/XHFd7meD7IJLjntrW+5EImeoteim1DkHQ+WjNOU6PeES0KZWZOlSD4UyBUV4
u9lI5AFi6Nc021ZOjdWljt+O2snWyFxUzkJKWheUkNwKIsS96wyWrqZtiDVpu5D/
h/6x/Du5kZxY5+iwHlW6ZrCFGyYemRrNxfrfoRCwxN8UAj58UG/74+Qmyl7QgYS9
HzAgRI8/cSGXBzY5Xa20p6D/1xDLy6YWvWdyCj/jwDueYP2vXU94i/KrTB42Amml
e03VZEe03Omx+6QcaD6BhU7AonGf1JtNByHe/hiNk2414Xc3F95elZFPhybp9R3U
nCK1SSC+2JxY3zvGGTdUp8nX3lzwy+7vgPaYM8cEJk6nYWkAKpOHk+yZJPy5Rfsa
LTWRtH/aMRmOGR+Ex+TozaBJIGEP3dn4rtIlZf3C/XaykRS7FT3dVgvrKA9cRqah
EP+yZn+qq5cuTl0RVprtRXIDugz500TstEvsuHcPLSade+576knTxMvBZcEcLEiD
ylimSb+HVpR8OnjLteOIVWZrANIzr67PM96nOdRmGnwUcS7+YgbPldTXPrgD13wn
OLJO2nK+NYi3mEj5dru1hOnGTqAdLCxvDzAeBlsLGC7cZtlXM1EU1F9O5ciOnMgR
Ij0OncFB0paJlDOU/J3/vgZjahNrwt+B7k0XWEbJrcZeZghAAygjZaxagPqjflbR
o8P2+KRnMAeU2+5UzAUtAGyF1WhYW3WY89PFJpHToqbnPTr2sYi9PbAu+GTyU4Fj
6U/pOi3VCJwA45kpcsY/gEZbuHas/e2Icva0o2L+bVZx5XFjMOvPkCE9BbiqfPbQ
96ozlbwOfEFQ1Wy/2Va16aO9za2Y77i3GTOWj8Lhm97ecKW3nNNMSYokg8ZzLMsu
sH/j+jzP9ibZ/ZM/eOlQyCRXWw/UASGek4fmXHBJ5LW0TPtp5iPV37LlNkWTH8dc
7HWiD40jLi3H0gMzzlTQuUnMi4BGF3U+JSyVJusono/5lQZRIX7nEgx9A/UQcXSB
b917xFBevGnUcGqq5pP1sX90nk8PNzX0BwYApl4mb8BH8Wuf3Nx6OqEMuaFL6bSH
eZeEGJYRS5Kd2tI1CuVoGyt7Obvd5jlDBtYn0dc6wV0/EVp3aE/jvl2GZGLGd0Mr
NdpTAoLHzdW8aQ0DrU9XNBTGyXaZl13pq8Rov0AWM8hyvrQvNgifa/BGLJVnwAwX
mYD2ZrWejczp30U4IKLpOALNBNWWGbP6gZDEoGJe5Ak5YWmb5VxFDmSJWGsEscJY
yuUeMTiNwadJnF5olX0sN/zzqGqAU8nB17embPyP73XG4gdYcvOHd7lwZ4YGsxkz
9cAIzEoCpjLpT1GIt8Z5LcSYeibTOllb9nOcwMd9fBPn6bI4Vq3EDvXB2FUwiShq
JSUdluWFrNJ/7P17tbg02i9afIB84DblDcqA2IHgumc80v6ZER4MUu8Sb6+sVOz8
bPd4kpUdKfH7mfOm+QP9cC8qfYTkHj+LG3LTfrgxSh1ZVa22lOap7vVlyqJB+Qtr
xbeqPNo86zs2CkU7oa8jajNpMrannMe+QK0VRv5x+RPRx0ji+264slH+A1qdfb8a
Fveubv94qxYEo6Uhi+4Kd/uDnqYZ1beJN/7StO3AZQArZF+bdYKYtyNsqWUpm4l/
IdbVRPJgSgrFMKu/VL1F35e8LSsCMpya1fa1eRfjSQ1cC3AAge8Ep1fs1T72+EqU
ERw64nTNrr9fx9V/gmKRXhyfXY4iqXRGCQS5faaBD9TD47R7LEtEnncJZbJg5EAQ
3AEzNVX1CvJSQp8M56CRb391fn8bJWOxFDgw4zXaz6cE8NF7ewTwSjrOU4iqFIxf
j9RGykmC1oD9HFGdo0IdIGv40baGlpI7SEXg1QDOvMdGlgDQmzsoTl/a+Dgu9fO0
9GnhUvD1qnlfKoK+foQjTIoJ3N2H0ZaV3X14l0oYA3zj5ejkyN/urTqlZAsCqCjn
xwKFVxzpJE5xpfuUT9ok0NP9HiuMFiQNd/1e6Id4EqK/y8o1bjdhxF3L2nw8IaPi
/sZId1aYEzR0iR8IlxN28mgY8HV2YinW3+3KvH8yTdr0q5DBaJdFt47eXDL2Y5OB
lIkkQlHYYodSgAulNZFJ24uONvGhWsgnk36O5d5pU/+Z72YDEYkO7ZIyK7ysb5c0
MEbkJfXqG+/1IntpnOlxqs7sFKhULX6O6QHg8p+wC+Sq0yBPc0USECAIpPMcjAsL
9y7Z5AedldtiUYmkemIz4u+gQaTYoLgQa5IC930Qwpy+hqI1kyrJyayOQWwRUpYo
ld3zPkrsXRPWCK/rnEZosn8M0KtNbfvAGdmjqlbJExTrUNR4UegpSa/8UL0TLRJQ
iEFF2Ko97UvN+ghvSwHn5kogNmeAlk5PB9vJo2V1kLc/lMor5qZB+RYk1cdsNDqq
UATzj7N7+cfcs93c0X+ClM/jI4Iz8vqCIPY0fWqcnOJx2UZRM4Yjej952g7hM8XT
OlnJVF3rTkuScQqQDnVMmV5np35e9NDMkgpFdqGbBUZtIvri1qN4+ZG2pKyEJpmy
lKRi/p0DIbb8T1bPgH7+wVSMu7wXsN2S3xV54sJaCv50b3ZyQ0/HeUSABviddBE1
IfN4kewnsr+byvk/kwAbrHxG8C7kBFpVh++FfTvj4uNgmp9AaGCYNfnnD232Uyi1
y/aNb+8afRzTaY5ySRCsIiKejfaQzwRPjDsyLtUkd6jYqBTHi/fghfzLkVtWENRD
jr9+Wto3jR81Aanl36wY3Xlt6t8YV0DGtNtisYXdPYH0Bs4QxF+8yaF1N/SE6S+7
9/oBNv56DMX/I8lmzU9kwiOpParefIkH9rP7QBcIUa1fDi8e/lf2um5n4RwX9IHG
vuEJapz0NZ24/YQAyl3GbMm+8GG4mQgT/Wo27lTBtATPkCc1KQ7E4F8hjYW4yQeM
++gv3ehZ4PX/SWm3/gXw6h3pkDFH7J2SQ6KW5O6W6dkATYzwGMyPI/QjPQlgzpL1
UQQO728uNssDT4zlgs0JHG9dff/m8pNYLRJbixdp7THswwP7lT7suZ5EBVv1oDYa
MxXXbRKeUN7YzWucwpPcf3CEFuvFcyIiKRarcIRj/xESxPTgH2xccdEf3rpcwJfp
yYoGkTJuHjPgeYPJygtHjNCzw3+fG80v5lTyk7gRsfTC6oYzy4kEaEv/VjQssWv/
V/LW5nF8jhrKkcpzBLiTcCrbEI0V12yPHgk5rIkHJw5gS8LWKfStPTD9ojo/kicc
EvsAiiSKpVBNOtdR/dg9SkYdZG5dEhlYSpAC19uZ60hWxAZJJxjpulvEjF1p0ocb
GCI4XbjS/L/nuwPOp5OumEfJuU1nDNpRwTEEUAw8P8wJN8z9itOfyLyIziRu/sS2
UbSI5F2jJbpl3J5kfM1D0Tdpz1vIdKW+54RzWeT5V0RkC6kedHwiq+ethhKnBbTA
QVicVVkhqUleOuyuQTy2trlk+vyp3pL6oIGYvQae0gqWKV5MT7nn46FN5lY16Bxi
2Kh2qcgc6dhbtHcrf8zvXZOrUmHDRRJRRmKcqbsPwGO7He5LOzh+1Bkeqaybszc5
gh128lhpAeYcAIaa2hFavtl4XjikiCtoA3ukErKsNURt/LV9V6D9s2MftZreTLOO
M9FLdcbXytjGH3WQg5RgX81Sy7+C4jx1jA/1MUYqkRrUNcAEnGEDqmfmvu9dVes6
y1rNBRNV75468Z+dnASEnEjInPnpkxePpi6qShKmECPLFSm960hqTyuOmXJZg2GD
XmbpHr4bka5mwd/vmpRp1gDrR1ISKqkMuuBV5/02Dh2PjpsWVLXHKOTFQhLQZdnG
wbQWFyQ8i936omv5dJJnNpr0BWdI/4xkWaca2nHwuMHey+jn96VTiqRfmzdmu0te
lMc9TU8ZsdSLlKf+oG+KJTA7SlpIEXl8TJh5UJ0jCjvqgTJW+aQ1fPqBjFZcMeJO
/xGILPpI9IhdoGCi+pPlXWq6jys4EPFKO4YnZauK44vNL49ZKHV3gvYrjrJ1VMbU
wF2fY4Uw1H/z83JiiOZPTp2eP81Hmc6wLbnmPn3PiZuWdRzFMGITIQy83YgqCQXU
BgkFJZSZj/RP0rqCFF8/JGK7uQka5jenSqBGbc5djU01KcdyGKjAcAxV8udyFNfz
N6n3XQC1fRoGvvBwx0llHK5awQqrBCwxr8kfbU/Cl02GFm9PtuNor8QCUBKXTlAu
qqs/ue//gfSfxwk1OZ+jBxeQA9uRQcryTT9P8r+NY5Qk0nze3IRTyPa1TKTaBUH4
8uB7IsvMrZfa2JoEEJS7B7sFOQyeYYkH5iL5MBLUgWAyHMZCBBqyahBTcAffQcN7
j8wmncoeyGd7HJ22XR+EKcMom56lDfsqbhO6GjcpM3BgGHKqDPcsc/H9Z+7y1uBT
ksPh3lczERR3FMIhOOagIYq0A0qhGPhRjwfloR0OU0t1I5PwZqAMAN+97bA4pF/j
I+Z4SNI3tpvfq/u+BFJEtjLay2A6WLrrXG7iYMYJ45CmACKAW17jAaxgg2w24T0N
zH82qim560fd1OrUQ+ji5AvKh0ahmzWeIMFoTEUnIEGmkPMFUANgzflo5u0sqvM/
/RE1N4MdfU/YEOrgHOX1nVpIlfqhCTtNSatmt/83PttLXUdhvJ3HuXN9C98JgDGe
LFoAWeuWwp7xiJcJLM5wAbcwo8UtrvdpBFxgG5Gmuul4KU26eNlZQga9eEXR2sw2
og/aHJWTmt8xlkeu0Yamdcb1txBF8UvKmRswKe41fEgfGOGJYsj3azlpu4b21mtp
6Oo0RUEFRSRVZ9b5iGFYKy3/LeLPUEPJUOwIOz0mncZakTYR4VF9lp3Q+UNdAbEF
aJK+0QfD312QB6wwCcF65BSL4jgA2P0YzlW4zgqvCOqvQDF9bTHGKXuxBn0qFEi4
sxdRizlkYE6PXxpGhF60lXC+/R9FMTdOMALdFH+8ifgENEBj2bT8dRds/dlOEBGx
84hidlGSJQwMUm38N+YF/bGegwyfFeHLN/vtHUxmwufvMzMsQlu5VsVdv907dVkr
1+8n8nWhiKcn9YodZouavZocC8bJIQio4tkHFqQSrHhZdoKyEM7I3WK5uGrX5uQa
QtLT+lgEWnLMg7tnrboUU36WeCQK99hPXJob6AZDR3HtPqHkrFVo2ihlBrT3Opv3
fUOoDGx5hhNMnv2r2/bQsdac2OKGCC2NN913zcRPhd3Yje0VizVDWp1bam93cJF0
lPMg1O6zHPmc7TKeNqDuP2t/DucOkZogIaYKiiqafJgvkLGIlfDTFZtf/8ELE7yN
wVDKyCAwB493ikmJvyn96IeCpnsy0pax1wErukqDOg3KMjiw/4EpLGY4K0U1Pdpz
9KR59gn2ccJ+7XmQbuWPQCPLCVVoPUM5pS4QO488CtJUjxV9gckERd4kXtLSLC2Z
/epWjmZo4/hzb+ALx1+MM1vy5JkRQ1LQSNVdkkdDeAIMM4RW5fQewYdwWxkhkVMN
YL4GcVkfLhVq7gpVk5qMcA1CbILpf1GOqv+2S2Umx4Ho7FPvf46tQUTosIqzBFP4
SOpsW74Hkkvl2my9xwyaZP4tjDdI4os85KR2RGWGoWVAApx1BW64bb51Ly0SJ+XQ
XTqeqq2JJGbypmr934qykvLkMgPyNrir3/R7l1DyBBYbYsRaBJtzoWN+8XsDuuWd
9UG+ESKdKeb5y2FL9QU8F/PAPPtnM22gPzGQk3DAaE3+dB5OtO14PaJWdyj4GJPj
g5chd+6tSjc3bhrse22T0eYDFR3JTWA6b6CjC6hoeTP2Oe4MHw6R1S986s8E4/Lh
Ueojd2cuVgBWojrwoVGrwt3p7PPCUzLT1Ze2Ya7CWcATMmbMHvXpB7e7lxz5b2Yf
xY2I08xg0igkAIqs8/Bs7xnBvfwT0+eu92+9TDySC0TG/dIXeaC3ESc3vBZIN0Ud
XuKKM7l41vDvZUnucQUTvG5aaiEGY9ULYg74uvxqqTm0GiUA02RHuRX+I0pgrM1l
aCYZ8Mz8hv/fpLnj95Ms9LqUBIesXfvTkYs29jFr+1RkuI9ZCNux/ElqbyTeJY0f
2+dLy8ZnwU+/rFzMz9Lrdzodyj/0sNV5hBUoD6xwfkfjg+ksB/l4h5h5iFbbr0kD
qfjy+vUGi4HQ3FHJYgAuKASO9kKoAUgIaAZqDtZEtOQFcXZ27591CeK41qy9S4E9
drMaZoxyXdtpR47/UGrPgvWByZSoXDNIkhSMwRqeD7jSxD+7R2mJ0EW8xK51UHjI
1wFsWDCx7AR0nPaSGDgrKBNW6oBYx34JWZS2e3KiTqSdrWXsq9K7mAd3nNlVa0DX
GeD+mNylr0F3tpk3w7ERZkQjc5wuyCOBe/hI2oHPtTLOqGROrJg5f1OYzfJamaGz
1QSosEF9Chu1TF3V1rmDBaDQHGQB2RMyR8ATgtUhg1wHCXs1vBpUm2KswN3kyiK6
FPl8xeg2dVZisrQi7ZFZyHn0SXMZ8NiWl/afJlUukBDghd3aM9SUPeFN47Y6IVtb
Jy6kCYTZcy7ACwJPckh4V+o9w85kwF6xcvYKPQaC5ZLC2vrEuvtJcI6nr/NLPT4t
jhMMGgj4q7r/8dMWnQm33kiptphCGRYCjJtaAhKp6ggV19BU4pCfpJyLhkvPgOWm
F/4dfnHMJGmfykqMwgCLY4hcFpKYrwyBpkkSgk1L8fmYSh53zq7hUrU4i5jCPAvk
CAJm+Cr9iI8AFmIVQ7HgLuYB9MmfvQSKm43xf4DP1Z0rPJJVzB60ECuml3QG3A4z
oZ1t7ZysAdD+S0/iZYdB+BsqwJIJqpMcmLE+biQPu7UhbEjwdYAm9fxJvoL7b+nd
5m9oIWWvKMPWRG7Om7Jl6qJKKD/UcfjMpRDWqW/sDmN5HZLKR2Rci7v01lj2ibC3
mDnxY/Fo0u4/dME6R/enGu6XrVgcoljVlBoNyASYyaSb3ZJ0RJmK+jF0bHI05ERS
VVubEWYKBAbnAdldUotmvVcwaDtXDLlc4/w7i83bF8NUFr9LaT8eBKmfVR/Vmc14
vmDrlGMS3GAVEs/8fA4eOjdvml4ulG3+CQEl9geLTh1nhcOVRRWaQuHJnV3wHlUk
42B+yJYJ9SpFjYplye0TSlWNwFKiJ0wJhPDkj5MSC+w9WAzlqhRhlb5H49UBlHHe
C5RK3nqdEvKPlu20ZVfwISgBxlgwTW0tUPowjzQXs6OvI/TX8zlRIyXU3E1vJ1VJ
icLWCXfUtuJtp16Dk+iof6HgzoKQwl8fELhhkkjFk7hBPR3LoA6Xc1UVi2+Kqi1V
lBt8S7qLlEy4c2OsQfG/QxV5VhdDQ4BRCJltd2pU/Z02GHciJLCNd5juUbA/IuDQ
PlMo1QPevcKFVHAM3zE5FfJB+jBOegryPWhPd6qayFQi9NTniPg5YVWarZAozWoO
W8rSgTwIYcGNuRzRsHQp5NgeTzp1Qp7xsm/xU7iEexPaYo8QaQjHnljJOGuInSyd
GdGMOCm7B6lITJ7RUlCRpdz3ZELC1Zb3Dn8+UjVh1h13nbh8P4V8tFy5rxGpjJTt
bEanvr2a7ndeYTK1NBjlvakFwdkOfJCPgGN1PvEj0G/InjUwbWZpUMPHSlsip7B0
bOOpgdq55LL0iADp+1dHIFrd+idOVwApHGeItqoqq6VZOTRS+SC1sH7IQB5V2Cpc
uIMvfUIP7WGIZdEzinsvJ8f2I/SSnzlO3yomXYQofwe+WB3VJEZ6STXImm65Apoc
QV/umAboUlLwWeWOTN/mIM78xCn5pDGFmLCFvU6y7lPXVF2reHBHALXcOUWhC2qa
u7BEpqg9Z2L4/OcNZDogCHvteBwH1+aeihFOYdCpYra1WIl91AOVMsy6K+3AmMeR
qXU47bQafkeTb51K1DEs0koFE9aNR7YqWe6xtH8xTHNsqyOl/YOAcnDLOJ+jn4Ss
a+ybQ+eewsj+MaB/YnLshNZE602qwPOZvfBOE+nsMfvJX0V5LkK/PLoBsXMPaf2T
J24qwae7RFuFWST8y+U61BDS9aHPNfs6ihNtEv3T9fdgV1eA+f2stqMjKLFHqhi1
bFxczaMzTXrFsu9pY4R6a53rZW09kuMNctRPRhiqnNHh1MaZQF8vsiYKtrhzRgGX
7ic/paWYhB55c61vNjXDDpUlRWR8NbVsP4Lebppn805uagjWLYlhKqIbfgOEfkAm
mlFAnhevL00L/SWbEhsGv0QxwXSmZwyLFnQ298En15PuRVZwWzRGE2FoTy0Ys0yP
Dc2L8GERKkEUe0FP1gAr3nVN3iFySjjLAzFRGBwcIFExDpdzA1FTin2i3CjrZBgD
wnsw2ZJ40gEVBfkkGL/wq1b9ub5tdbVdcmpraNa4NQ95seqF8DoYEEJtwgfbXRgA
hX/2HI+nf3kwUXZW2P7eUl0AXipvSkAtm1PxkBrGgFmU/ZfbVnZtCvxhWYnFQQxF
92YQf2IDtyRd2zt+fdimgfCaK46VJcugYHUKDbU9On0Kyn71dON902BFyLfiodPO
NjhCoZ6zHiYVYUxQ4xLthAuVx/yZmEcdV1GIrezO1KK1oNZMXvRFYcduFgOQt2Zf
fzXggEi1wC0NLZo0KbewRDbxlne248Aiqdl1DrUSLeQBwTklqa2aExO7XbD01tce
U1DL/GcSGFNda/J7afkI13VE9hEj6O/PEIRPyXApohNafdf1eY+bOabITAU8vj+e
JCufABTa0YZPqkudd7zeS5wgzTulApTnXWy7vNkxUg1WP/oJXGr804KHSGPpiKXf
5IqeiFEaQNU1QmkxCTBjvTls41d5LsIQdWc9XnUOOjo52Gr00jNVo97kxVslg/dP
xMDuunEAUNGqz0YfzlRlXDhm+zeArNFwkJaq23N/lpAjVFPEMPACCUmbLyMYZwQY
/HeXrvMr/YYkRb0Rwjx8FhpkUXJ/qLeSrSG3ehk15qMAsuomLM4cMEjEnPkKL1K4
K86brgwRcA4fUKQoEUGC5k3sgvGh9JUYFJPe2OJ8PKNVPSz0ss3tdptRMbwKen3f
OB5p1Niz+fW2svl/wnqFrwFJFfYiGActtIf0DAp5a40AjYko1HsAyk+5ep4aZKxK
oxLqM76Jd1j7L1HCGevgoSGp5xbayYK6MbUkX6H2/x+/Rue85XIA2VOv+y+HdE06
AjiylvcI+HVwmQtUp+usfiJztjgoFqEi6qgHhS4G7knuPaHqXgJv30RcdYpKC4/V
rWYHF6m85kvIo4NkqDnvshIzbVG19Bn9pe+F2Y9bWBOwJiUU0hn37lERSQaNJMFk
z4HOP/9PNXgRaq+BdIqg/HLG2u4AGMUvU9ZtmBoKaLVt8d1ZH1uUqDUUguIgOcAV
9USgbhX+4FFQG9bDEbSSOInsEFPmbt+LXJuTvvg47CkuyspfNlD6isocwLj6LWbK
eXT1L/Vm0LcUcJt8Xyc8qWE+uQeL2o2xvSHFt16A1mCh+vUTfPJNQ6XTvG1bZmm0
OiZHZbYx+52p5h2cFTcWt6UR3Cfii/9nUB3qv1L8pQ/LWghcm/CcilEfrLDGAKcK
osMZSlz+ibBsz+d9KBpfdS8hGxgnQFZqn+evW6PauuHAtfw0HcUo5/9rq7UKJnvp
3t8sVo/mP+svfhDa3Dr1OccBiWqKWmRF+tDL6pAAXW1KFlL2o2LXYnOWGTSPm+Dj
D4X9lAGQDzQTwogXXS0WAtaBzCTu6gzoS9kPwcaJjPMo0m3qmzJI8421d+eYEGoW
/bnfk+98NPqQbyh/YJbRD2Ye4M3EwJoC+f4CU2PFYJWKLA1jDJBomFH753ZaVwgO
wBwQCjumUEy5ITbm4j/C8xYvBFVBt1LyeINmQiB4A8Ip0r+bNKO0Tr43GAJMcH4d
lc3MAnCQAAMDOpfcp6A1yC16nH9g9c1esS2nvncNEp+ZClgin5Pm+G8XLdd8doep
Yumt2aY33eJGf2wa+eg43Habo+4NIkPNJHXqhoLL/W9r36txjKcqIJ85iVrxS9sh
fd/VE+aX4maKWrH+R2yXCkSFyJw48cvyYXvRkLuHereAQH5QwlWBYKXCfLjGG+fS
TH6nl1vPblnlVqGQ+icY89gvsz9jx2TE0Pe/3qERP2C8bzbQSdf3Gq/r2CPYLwa6
YjLKU2OrI1mpxBZZQIgmw394A21BEfA0+5VSWQHomsEtAuQQrL5NwjdQveqY6sY2
aAS0NJ9/1LBplEy7qoEYWiayfpssZDhcSjLYIctNMYhNP6kNkCdnex0c8M/y2BPl
ngYzOqN8eSqrH8zTvF8i/c5m2Uvr+LRVUz4FRy+Zy4PN3uu0rFTsBJ8QWlJzDU1u
rsNfuTPvP4twQyYskPBRpxCHXR7Tt/kKZy6v6hI5UgAi6bpK55cavWQp8W9czqBq
uy+t4q7UthG8C65ajd6CJcUkd8EWh4oHHHK8ITw217940UQQ2HcmQHb5cJpliow/
bYaZiyXUBkLmZ5vQgp7gkm2iI6XMntSPSan4lwWVi7gk/se91ftcEKSE86EcJyg4
D0ciD280nqbdcViRSABgu+RHu+XGiq77/gXFFvrPIQEczUuC1ZmNu80r9/zjk8ag
IlL+sxnLwOzENpQLAZrv5YrV857aRKotDkIGSHuPu8LSvUySMXxW3oFUBEQyVsKg
SZu8nn5WRHFTIBGgK+wa2nvHQ7XzUmUOFBSYsFr+KArjmo8JALLVFQDCMZiULkSe
oVxmkNt2kRsE8H+iKUbLapGhrEZnIcmQrVvbIgAtDhzrOAIjB9Epl7TsgKw0Yqux
yUmJyXIxx5FGfZds5XUk/XfHV5PzaA22BK75TNlh80+S62qfZHBDGOFEquIeFzG1
DU9ch2fODjqGtJ/p94+WF4Pv4J7ZfT3GeCBb4sqQKl+I1CtmGxL5ti0JDQ0oT5RJ
hKNKGt684WwJ8h/YPUPieVHCkkFceqoXxkxaD6MMtAkDaZYRkVoHtKFxZ17Mefoz
ZpB2GT+eYaydQkFEqPShs/DjhsbROKrQOXE8AK91oApkuh0993psoVTBX5YoGfEL
dGFjV+aZsjT684G/0bbPdHWN6h5W1iDSqD42Tjf+Q2Ax8s6171vepxPDTXD/Q5Ia
VIPYBzUbeUstkjz2H6jmWcbVvKD2Z/IsPI1BNM5mY3k/fWY2kFNjEWy4zrMTR0/o
mPL4/VZdlaJq+DumKO/0ADL9LunQYQmPkqvi+JmtkXmY8GFykTvBkeVplSSz3POW
A3jIOe+XucTKR9omrcBHPIIA9Y+j0AQ8FMNkPouCBlmZwfxuwTJjv2ET7B1UTNcU
N/YWIpN/JNuZbP6oxgIN+SxvlUN49+9yE2lX3X0Vm46O/Gp7EzhcRB4bwJObv9/e
18pkjXKVHKY+6gc+gfLzWOwHr/vHTNMI1xWDCin8R9wv43zLZsJsmsOFkE///zhr
HrJpWOa5O9xaAdM5ryVygUoLijc1ezSjfRfpc9yX0SqamQ/f3cZ7fd6VAC4mybod
obIXHmll+8n44mwED9QWTk3qhLSKeD133HPpkVzpvnTrBZ6LcsWx/8Dn7rT7g+IF
ORUIpMcnjre0TIxvGuGrp1nYOF3fbOuuZslhZ+MBsq9fHynHN94iKDdTHWgAdPpQ
Mnmw9sSAHWHUMd/Y1d2l2Ahrg+v9PSG8xchp6e4cgo4TNDFA8bNeoYTacI8ObCg1
6Jj3Uk6IlzLLUKJtWBKMM0jh4HccwuwmXbo94bvheyaACFUucHDH3eGfg2PL4sYA
2ha9kR/6zai/XzZj1oID7dJh9RP0/dhSM3cUNsrhkCiaL9bjwhkuI81WK0WjjxN6
TYy1IaKCBnkq9F0l3sNYNxtJsidT8ZpytFRTP3/pb2vnTmbSsCIrTUulbDlG6HjJ
zuvko0hVjJ5Cc8m+D6UpQ0uiJsQ7cIIeBvKvmRLYeN/9IobEeMRywqITl525tiHV
R+wTDrCeBIkanD6mEpoL8DHLc98nJy4tX7mbZqITSFboZQD5w/23cni48V7tvXeP
QZ2SJg75YTDoJowEfS5nq2DQrRja4VsKCd6sdrlhSS3wAOsJ9h4W26ZzxY9gx8DU
s3gR4m2M97MAKHp4CEX+BO7DcC6pjueFc1FkNhEQEgxGjMmGI7mIJJOdxX9tImca
8X9NO+5BGLXBSfN2YmfcPd2Ande+M8Sgpi+VC40xN7dm95L8v7+zrqv8IsE4mWcA
4VswlGL6bfWi2cg+xjjLs3oziatUlrmKKWNBm0MLfjJb0q9AOQzRfoDAwa8jGwrV
w8Vr8fPuzKrCllL2e363rooBHymNPeAXxu2ut8OMo7NeuZ8Qgonypor1u55rNcjm
PxfBzSfBQzs4SYrP4THHx86W9eTPDRWJD4cljBBYgH2Pl4g05xinlRCKKngOjKN6
fUY08+35rA+PRjYHAeCXFm+xz2sjHqZH72B80pn/U580imqt/0R9nYHvEoVlz+Fp
eAP3NbmNAymEJ+NhxteVYOjEz7NSJqDEeK65RODVYZL72Ze8h15J3XOh1zH2xijQ
axlukMDaAVwHXqxvctl/Y3cSP1xBPfdXkvAWMbZEDdnUBqbEJgyDgK0TnBluxc2q
nZJeW3RUUzx2kg4FdY9Zm7EIHMAbZ7pn/YEn3UEQJMMWh9CYt+oX7LNP2NRcTaEV
JPtxiCdCQB1YsAlccSilDlBCX11xmcEnuUlFZwNWLQYeG6OWMbCKbjcEQGK8gfwr
wX3UVgxqV0DV77urB40aVKSv29H4m7Vaj2Lpmg9DbTG4hcxmGC5qtuKDMOQ75xDg
R1CsISztZS4VP8zoMKdrH68fa1slRNyKHAY31s2LwM4nkSIGwu+5MQABLsN7xb8t
v+sYGi2OaMtMcXdVFq2ae7EXdydgBrp8+5D4sYEfojL35oatkQQEwqqCvMEfrlQ0
9lpqHkf3MlA+XcB7pRb2k+5vh5/S/znQ0oTIDgcQmQLHtbXH+AgkDXDB4Rq7QSNF
I64HybkEiX6WePtMCAJyk0urLjv53HGPUUpCDMAvpATXu9EsgciHP+AwjQfZDxSR
aIwT5S+teLUF7jvU9deuFrgjhG4zoGzU7y/IAaLmT5JRZZlVZGzeF8sp9m7ELDv1
cFmPvjrs03OKWqdxPZ9zfu5MeZA2G3DlUJAmiHHtv6XgHj26VDf1vrnU+LIylvA7
Wz5G802kBUw5HJBlIigcmrQUCjprcxmZLOt/l92n2tJF1r93kteZDLyCaklOymq9
mPf1qVG3rDFNFu571kcG81QPNj8pCkOpA4l/BvWqNfojz+nMXFpaTG4+pTHoIhEk
zWOwkJnOkJcuDHeDCYxuISk6loE21Xwigb3qa2IDBF9EVFaK9Ig7BxKiXc6XurAo
7HOknbAsjcwchWeFkUWPuS9mhTivauqpZXIo5EXC6IQSuMBMf/zLOCrhLuk5FkFW
jdXNVlAbQc1VgRdWe1QOv5L8zAVWKpBbwB3pot+ilqpDbeXCeusmYxpn5AvD/XpJ
XHnSF2X32LQKNNNLQc3uYjAytfqf2HeV56kHeFdcqrl421BZU6xJLtmdbM0DpUPd
LIUQT9uwhrP0Jcn3qYeb0otIsqfqT6IDPfLaGhVVrZvAo1U6yfecu7L689Cb4Vbu
5BywdopjiEg8PC/Qv36K0gvxT8zHIRBvD5K0XDx2ro8P0d4KHEYbDJscpW2nvsPj
6OdFieWUGlHq+g5ZqBM+PwZ05udWmOdaga+eJw7DVxNL4YeAczw90bb99n+Hv/hs
GpSoJKg1Rup4f6WY3Thdn3TU1QWsd4oLLZCVDmCPZMcG9dlXcD4NSQQN+iQiv4Pv
zwnLS2WlnEG2Mj0C7AIuTY8cJQB3pqgkKzyISTGW82OwpayWUxUJjAJlym7fsm9c
Hy6RfkYOhFZpuw4eu4yK+N8WnsXuQV+ZA5JAEbREh2GKY2vzCqvq4KOzoLpcUuBh
ElJDG8CRHtefbUrq9yscCuKY3+hmAIh2aFfA5D8GFBpnEcyr5IqqonpJo9o11QY3
vM8qEcT0/ERbJdJelcUCAnSFlwK3ZRQ203oJdlrDUPkKIn+6RHKm/A0QwfoKaP88
QbHTXmcR9TgVpnP5hQs0t9pu3jhNIYrcJp/SsOo8PmhxNDQol8pjS+lWfuM8KXai
XGwHUyAi4jietLoitAjOhYfzsBX182AXDbhQhrIWv7JEZlnn1FnWOFyQvWn4/LWW
VvBVTRrpqrTOQvu8BkYDycKq2AhDo2ds7Pa8b106asYNARKYFIswRayGUwEmY46t
RTbIptb0lYHSr2xPstIYYA80/7NQyswBFOb7ZRhNJ2/RXxDefwy+HtlsRLM6nGnu
WHoolRheU/ST7gq/SvhogiNPBV+0wHTLud1r7rZH/rT6a8nUo+UN65PwtJRNB3lL
+jkxpQACPfueb4o8riBg3M+EA20NDlzUMRpmyILqdq/9mPO/SBGfnKodjsBdhQ/s
L/108U9ZYw+xkOpxW2sw0znQ+xDQtpB0RRnNJBpR6k9v6CmlMBpegsOCzEg5Q968
AMM+z17Pei0so4ZhnaX1zyrHEdwAJm6NtdUvKcN7Ca56CeLv1QaKsHRzZkDgviW5
Yi32CYtfQjjZipqtfM3b2CnzoOumS3CmH5uoc+w0LBdQT6KaVS/mqTO0K8KhmcXB
phOds5CnWezMSIW1WLOU3xV8Uk8l3LIN5TbzzMaYSB8e9xGYo70jG+jUlVwlv12N
GQxJsTMT+Wf9rr3/OjElNf5LMlVFlKEy0z5n3cK9YJ5iFm02SeqcdrlEoEt2JpoT
1qKVJjqZ/bab56pO3MzigD2SOYAgqzBizalY9Hzum4C68YjsPIiuNHkc2kOB+eQw
sbMi0m4gg4tTYGOfOhtYoZkigb3rxvcDcN992LPZlh2s90m8VMeXzdqNMQ4AKfiA
fA9x9V89WSC/UtozJkAtnBlWtwCIaOQYoBHIcQ9T5HYJguOt1l8dajha44D3TcIc
ieIsyGdc6kQ7O7GiXDUPjoK9hvjI8ix/T9A47yVMRbh3NkHML0IlmbpLIFuB1OhG
PqmlBWkq8qCDZF1VibzIXm+ysbMVpglNxyNwo2RYRWyTtxVqMhwDElVT7v8+TCeX
AAPLWlWwc3pOw3mU8euJWtQJhgz7Yp2Tjv2Zhzno6+tDKnjkIG3B4pKrlXnSkpOH
gSxA1jv9AJXHDWLL6AU/2HYdoZagU7GUq8X2K3N4iMeB6TRbR8Mi3NjGBzp08ksJ
t8PrRxbGDzn+Ivucmu3ANqCgaaqwhxIoe9Q3A6+0Zl3dZ1DjgqYnd1sVlgzkBAKp
KZKoHi4E/wvKShUb7YgVV7Y1p+BBPGlysoSs2OT+WhHIDDLzwhNRxK/Nd3neuSM9
kuzhysDGDjeM5vcA56Zuu1cm9XER1G79xAx4Rw4+TYmvBuNTEgKHgJXwPhYD7XmB
KrTYUGF2sFB1pEEBnqbSy6kCCk/ifpbSFrhpiFmS3twvqQcQUIvlKUzmSMWGhVpX
IcDJvmprAl2BctqVRp0avG5bPuMb7ZSRRFvUogTKyL9Kdmhznon9cqc47xoG6q/E
RKmom735WpO4IiFoO0G/p9aCLgSqW7VaDGO8/ok2rkTCpk5d7B8teoa5lvaMsuoH
xDngcTAE6Cr4xeYpVZRkCspdAnFn/AbGgLiJbm+TnEQgx2mvbWJCbrPPP675/mzg
+1mkC7OSM2MAhHO1kC1qWANBC6guZ5lqhbbz0hS8FTEYO9mGFK2D8RLBhCv/b9qb
Z7tZm+nAWJV12PMNFMrfyOS+vQqlf7FODEp+FgNTT/VxnWdv+VzQwCzM9daB+H+9
qhaVx0d+59NSxxgphK04kwozDUnQH5RrhReT9RMEtSgEpSjm6rNp2csIcL/+K7UT
RaL3gMLGLZkh0TajewFo8jplKZ8Fo+uq6pCKJUT78r7luahzOwsSBbrL7iNgizrg
1GypoldpTmujJw8ZthhMfTscsTNPIhPIQ9U1wNAm0tQ3SDNLhI5otHPBRIDSX/pX
tJpvCK49LuOSjsHOSSiFJSlLBxhpwoWb/NKxLOYoMgEe7c17nt7B7dfiXmXLh1Pb
UO6csnp/LYDfY5FzIfRdz8z93vyE/wQgqgIsuE9Qk/fHwLFJrBg65UnoC6KxQMHa
eWaiA63ERjQk5XiugLxL7yUYt2cLCRMOsi3VptMMNfz4bkkKT+q+ngX0yx6F863b
lbUYudxK7SBkaLxd33nc9cFcDHfySytvnLYlZ5VKBhtYE33ChxwDKU3zit26oKpc
8D26ElNwXHiiORliYC3QOu6tc2AzzXSJY587GiYF97j26PNkWA+8445JUhKlI3Lf
ndVnp/EzSCqddKKRO+aIQQ4HnXfLfaaTgdayCh87xcojTY4/Qs0qWzJ8WKLWHkHK
iN+ai9Y5HzT/lJlr1TwrqKNRbaeGkZ6oRljYaGt1SrX2rWsKZqKp78LFceuY20Cf
wqRvrKbISe38M58yCyZdPiUbitwJFnDkBv+bnzq14jE1aFLsK1xV/kIlAJ8iJqXm
wejTa9Zmz4U/97vz8fUPdd8QV7XlY4Txm8VOlstNoUr+wfrwp0jxm3HG9zpn5VdD
JtvjDXLmdcanN8cBJ1P2Pdduh4deOpd7bYGL3z4D5nzfkfdHq6ZOTG4LKIY/v/Qf
I3dvaZAE5+tqsiPHrwP3N3kWfPWZZY9mAEKoSGkjKtL44N0egArsYeIy130eRcB5
K7rXQay5iMOZeRD66wFeHgcItIbWia1+LKyHH1Wi7q1JxxwO8hzja7egFq8hC4Ep
fv8mcOCI6Aa6aw3hGKTQOepAuS5rAdcCAUHjG4gZr/SiEDdtenCTrApB6Svu/325
HPgbH0b6Ccwf4gxuvzBh67oUUaJVXSjFPM1NUnMkqQ6ginOwp4wN4n6ci/GFx4VU
eqD7tt72F8DFICG3m4THwLDw47n4srPdQS8hW59vHQjaIftE+6oJSmPitX3PEyXR
/JLyxF21Hks7N7pZgJmhOwbXLzKfHCz1hEMI5vSAAsIz65SYOGfRp+F22QMaLLzf
zcFCsD1Dfxzg9kZyqmS5ObMbQWlDSmMbmhoA8jnqZJp9MZtjGQF+EdnZdhHHDXY2
0eMPPhbxOPyXagPqq2jFFHdD+PJAN1vYxcqR3K4EN1C8qChiEZcf1SwSUp4VD4lH
wOCqW9FRed9fBjyIaJ7jSNxbG2WN7ScwUhbr01Y5EWOvnYX86B0bZcTGQatw8XfL
zPkfUGd02SEg4DkqwFGBd/J++tT7ICEoIs4C0S8nUjoZA+mzswuPUZahSJiq8ntG
vC+s+TTRvcA6voiQc9RlbVWX8RA/XSZaGAP/C7iBWD4t5r1VDs1eGIUc0i2IgXh9
csCIr9hMQa6p/2N24FtZy1ulhoKD68g9w+F5fs6IJrU/74yOwJ/E32lahx23wBX2
YVeRbGnXZiSyjy9mEUXzUAcFEiAxmCk4Y5yqwgMR/FZCgmypl0B3X1kfZANmS3hE
WQn5CjFT4iEf194TieJRIzvOyUJ+xtcU3EhkTT3KgN1vABpbUnGWB3rxI1QSMWOi
H8cDiZX8xOBykQBF+tIqd+w73K4dRxqgWo+Or8YeVWgwXXBB45Pi1iw1hrsmXY/E
M4Ni/yZB8Zx5bm+n5s5Qzad54L9Dk0O9rDvtEJWui7AHdeafQp6ude5yN/ApcAeg
DfHGhlvvnXb+d1E/VO2LKIn2zbw4VI1k8GMs4xTD/8uJPTzQlaMORzqdc4KLfeRP
q5FM7Kf/klUlecIciPiJS6p/Hwa94ZDXq+PLy2FqurB+T/LwvQNKTuvrUrgVuHtH
vv6g6ULMHQoI2U6gi/NY4SR14ZyP/HpDeAp+ek+vgHuSejfT02csHFtPcLTYvPRc
1OXc41dacwcaTLJUMy7CMh3YA6SAOshQYCPuamioZnOqCadjr19LCvpCrKKXsf+o
EpAl/tpYG/ALalCYe9zVmXbe2WXhqgO9xqyWrTIaF1HzLoZdgR6Lcd+zXVVxLwu7
QX7PxRGemhev/zxm1EWEtLWrvc0RNaIGrDdALOOdds9hOFo/LL3T5RVKL6Sqf69o
R3mD05l6dBe2Oyw8BNSD6H+mFWQaOc1F/lhGqkgZa4ZlaPkyDiCczkTEQsMBfBUM
GKi3O2Z8ghudSMxK4atmlPkke2gk6g0XqiIdmO5oscc5bZQQ6vajWuHQZC6aVIux
/HHQMDCHiLEqc01IhuVAWJPS7wD896Hfv363meMfc9QBK2gpdjKuvVOmVGcXf6tu
PyOSL8Hf5kUDs1qXYWN3nMwFOUyf7MzgyCf3Ukzr7ywCMHcxEEuXtr0/P31zEJPp
3GOdXELKZTuLB7mdpOQXiWS0s9VdY0iaSENTCp6ROHr/JVzKtV7Dt1lwFnSRmQkX
uqEW7GGLbNsWDshdm+tlq+qioWCStLxsMjKE4Kpo1B5YH7IK19niDHSnTmqMeArt
Ml5TKGxQjWboQuKpL4W/v5ZlW54jgoHCbsetB78OipFjrZSMkUpSyZHc1Y44/USJ
uqzQ1M297n+eFXAXoSC8wr0TQmMYYOG8lcTVSaQOELmn4A7XDe6hWJ00kny6iXUg
C5rF4BHtVZNZpYEcqj8e6pLQj2aR1tPnQRF/GZU48BtbnicK2UQu4VRyvsostHwA
6Pmthc5FsGUyY8ktZDUB05MAD+bFeWURvhM//EpaKyyx0mqDCj85F3gIWBenevcn
wnv1xAEP2F8kAtFjYKnVqLLxBJ8ysEgl3dUIAIXoPj4n+k7Koi/dFZ3hxno/arex
jpObO+DEQIowFdwglMIvSPFH7vhxDzInoSiuD0+dDLUTgOiofMdqOWSUd0imccVu
O/F54ZdjmhLXkIZX9T9EdD7hxpWp7DcKZgK5PqibSXwZUSwi1fWMdr3lqgfSwg03
UOiRrHPoNsG499D8suE+lCqnPkAGDy5g2n3K1X6lk/mbqfPusmugizIBvTDVqKU8
nHsS40qPY5uaCcHrSgUEygIs0VUOKSMWf7Q7EA3nuxKq2aJfsLKTtL4WUZHbRaOD
WjWoMS/aqbYALuJIWrl4AxDE4Zpi3V8tz7utAiC5LcwPv6879zE3PtsBoysFdW58
35n0y+OtieAACC4FLNFXzi0BIR13rwgYB4nTNesxq7wJeC7sSpcGPBtB5J9qhqOE
FdBUb9ZUPgjtwDrILr4TnglQr14v8YWyfM7q6gYq/UqSEIkaxEsjrURINiTJYt+G
fFVBUM9mKQSsUYBgVucHg7xKfzIsITUQWB7pr8BMk1sAOlovR08pGMBJcCKgoPA4
00dnim1U+7Sula0WGudcWzgS4V0E1k+c/k+vUoXEwPIMpTgJxinjMZ1focXAXDN8
vLT4i4c9fYS1qCDxNzOzEqVm7MvBsbyChEP5lgOfXuW/5Jvf7G7mOMz2hiW24kBT
VmzSgWTV1UG0ScuIz4Y3l7LwpPKutm8xDroWDY8/ZyFCcUHbhibdyrtAU3JInlHB
qzc1+/ucm+l6L8eKyRwIDFLY4Kv0Za9+wnhFJRIqzh6/orawgNhwE2Zxrdi0aIFf
2p+sX5TkioXPD8WUZcDwJGa80iAuaWFo0srhJ0OEa34ApWNEgy+Pxd4mQ6Doal8C
dTRyrvF5tzQF7cwBmwZoHFfvUd8ipmWGcoGVcRkFPajQ7xg7RrIhJpNcSlpCKaFc
+y0X9cMUv1s+saCo6h2N11bKOqLeM/zd/4XSP9Uj8ln5S2V9THm4RlMQpjCgDWtA
4vToZ7KIsrDZgBSSmfB6kxYFdUPwZ6YWHd501sm+q4dx0tgBazKPVRg8duDeAASd
QzrtMYQeBVx0O43ASPYid95cCElUqyfkkpoPxNg8FZjgqkqypMESGjiFRrHiDwvD
1GqVM9Fmx7lNsjF2SH9I5+tsnqia6DbSFm94NDY02pY9mFNgkccWvU+j/aFY5Ajc
QHBjghM6zGdl8SZknWsbluurMf71wcFiYYYxzbGsJ3QpUcMJSaP3isEmRzLM0B+u
rpwnzY6Nc44h9EbpyAwm5UgnEzpjclvxKNwpYvNMwe0q/kH21wxKrmweyB1BMNFp
IvmLi9Ec+iywaON5YB5iZw289ozjWBnFRXsotuJcanHnaanM7kCO5YjLOjobQvzz
sskPfPeAfRrD3h1Ppsyd9GVajsuX2hwFrzkuv9sjC2aIhl+XDCm+3q8SrnUd50jI
SRTscj259FMiJUPD22p9/6KJBjoDEvjcKmxfaLph+z9L17naeWcHK4CMSTFg7P3I
HCXpocO+dfvTihjI676eCQR26RNhfjr5VWaiHrp1N70Lk69GMVPee6/y6uFc3fwC
jDnYjB2Nmt/MlOB+GCUQPl/lHhGQ/ASv0NJ2KEVxBaq/pHuQwJvlphrdi8koQqBo
mRxQuOFcaJCo4WqweabqtsGwqem93y108PMSPGkuCdgOOaN1WjSBHOd58ePXeeSF
H9hnLTAtmEhMld37GB+k3iUKkWm91uDB90W4PC1/lnIe/emtcDxtXBFQstlwm12m
HohG7QiLFoTbuaNVGj87WMcaZBh9WbBN9LSItZ2MQl396pQxWZihKLDUjwLlvl2s
MMf9dXL1gpp78eXeefmhlQZsHU++Wd18MKbpN6vAy8ejcX5XJQVIOVsKV5DZyy7M
O60CKxZ6RF+fYAnwl++LWGwsd/VitJKcN6BufVFInODd7ju14ViGtEvtKsSQ09vp
RBGgBGq7jdJW/+ZcRpzf465KGdxhOpfKNACGQRxUqGA+jtgVwP01ZsrAFOTWTKtJ
rocGxNqhJbNkUhnrWV83BA4p87sNmmkna7Utg8zXNUX4XDrmID2o9B1KFXL6ZpHp
MwSWHuEDZT0zxI2UHM/z1j0EDpoQzFgWEsakJfXKRkeS2iQ6Lq4fjmYTe9m43HAo
Fekyf5WKXkCd9erPG4bc3ceh1GRBKT5VG4yPxTg+GmpHgk7TFl4q8gV3PLaUctuM
BWju+XGHLkgX82OQJ05Do1rykD7I9SvufkT7YPtI8qDLmcp11mhVQTKRtYuZM+yb
sJnScRdHCqFDjZWfr/xT5XHgBoCvXnW6NvgYKFI4TeB0z+wAg47WolHQ9kGk6sfR
MLnMfwN+SSqLgPUaVHkbTM3WC/u+0S9sAH7gGSGhar7b8XrP2UjQkyHWu0s+Ee/F
or4RmADHQ2Gf/PpG8vMoWJHoRh0/jXrn+2VjlZM2OBWLN3chZb9cFAjt/+li0iX3
lLcTJVFYY4gPdY4BOqsWGZ5V3uDW0Ij0vnR4KpncLquGAFNlkoQhkIZL/+O0CwFy
0x2P0CW89U93OpItLZcyhQABKG0WZhHGCBUEgZ8gRSCHepbQrOByjyIK545DjJ8M
MI1FYayJZ5ciGBxDXPhIlnMqDTfRlAoJ9eo6TzpO2NSxRAn8fIVGxz9Y4qitO3xC
lVbolh3n5qIpO49iSRB5s8A9UXe30vzptOg4cf7UUhLkyM5NJXZtwcDtv20fRJIS
ztPka0TupNjR9rYLdIy7ugk+bImshYmn1dXZ6c0r9ulmlSRmbBNxQYxDkW/4SOnP
ED+JUZUdSrnISWiCNdgYwNvBhTNIWpsloGvNDA6ViofzAfuYE0ktXRRz4+F3+6De
XafNFvUZY8yTuIVBGW4AkKZGIbX3NL0WjgSh5muUJfrPHAmcVowS5CT0m3nruVY+
M3hQdsyeCBiwJ48ckpz0pPfqPAE1Vukv3jCk8Nu9ayg/sMIP2MgcPo6rWDvwTtm/
D7gnAPP97ZZG0f2T9o2KQfDDxsMX2bHRcVaApHif+HMVK2pw8gNHbmto08yQbsTZ
H3tCdOQn8/uBmmy+RwPNnwc93T80Txt3CT1AryVr0fpJSuWv1/qk1MTny86R/6JX
JkXUX9XO42SDOrV5C5rQp7XsQmvYSsEqsPpiFMPISpplaHUFLVXg7jvLjhEcg/b+
mC1ZWcOxDapFXUpD5F/TQ39lMWaOL53tS7Ok9ho5im+MjTVAQF6QNMD0hVS8wZhB
4PPxIRPkNrJh2RaKkLJbWOkGoSgGphqdj5GLOHCHMqfjOe86uiwBAcIdIKvZKYGx
jekkvuNlM/EDOzS4hQ+ypYZ6Deu6o7zLm580roCJjZkRVHDXSWtWhY64cgYDOMrC
+31nlNnY011OTdxTEiCkRf7RZYY+dFRTLVaWeH7tC9s/BWaxHc3jTlGKumGik1W8
jBifAiPCqZz2NYW2sHasD+mYbBtgUSqZIeJqXdVVUFRrUiFkE1JuAj0oQzkHCmQU
DEWbx5CUVIP3f3dEQKjIUqdC9cz1NUJ5Nx+QADl8XAx4OrX4TCqIifzyEkvTEXkN
k2wgCmsBYZZDlT99nJMQOumwrE0A3w1wLHzCiyaNPldAxCKbAx8piMoie5d8hHK0
bnSRXKyGuO+u3oIRAPDv1blGyuRGvzvs6Gz3eLuykTDVLU/2ZSqw9JFwvzllm0jt
sDbBb1Ng3SLrXpz2O/WCzx5zk7LlIgpj1KvxNkIIBlyp2TdxZ3VmnFu9K9koo+jv
a7lMi8oH7vpwOeB6ui0IB1UopoZzhRtvSOyQGXkIXrOqZ3+QLOBJqsNHVjHxZrLZ
srTy4EgCX8WjCiHAo+D6yriKbbnisZZ/Wqqddr4pbn4SE9VcuR2I4kBr+cDsKtUW
D+xZK+TenzQ8755UkiQc6ti20iHcH5tVkC/nXAEMmMwjRhb2OccchPLj89/Xzbs1
OY83hSZxnZ5Ubfsu6tJczcr351Xc3yBH1RpA88k3gB4FehxAjHutE0FIjywO1YXj
W8MUattRd3GPrRMC6w/gmREB/hprTKMu5Jvw4VjiDW0I/qawO6ShT/TVccOq4nvT
FWLBB7p4sZChlKgUOLDGHHW1Z1X4pwzzQv91f4ASxFS/p1Ju7EDswrlA8mbed9Y0
YKwMuqwu53d5Kk4Zmmga/dhIdw0Qm2kVR8XAgvioYfKd9v/ecUZcTbxG0l6zWgeM
+OO63359EprvECTOUwsTXg45z02IR28m+M6Cl2XUPVSK9mtdmNlK9diKk9SH8lyX
Ml5OmStmeNsbRXBqYXYQn5C32TKKeNiU2F2G65NbFwMGuB0OpGi7VOv8dFDefDe2
VLb9/QiBsBJTNpzDEHGZYoZui/EEvkMk1b8CIXrhZWsT4escS97v54bhLfPzH0MB
Wibw5ud2LxovUlGqnD4v8p/FmuCTWvCUPJWqqOZUcFAJKd2un2VHdpheApA9t4lk
34CNEXPm4ASdXNQlaPLkDdyuScIpkx22YghnRsb/Rl8b/hUahSZHtGpgf4wf6TpT
tXx7N0BFc5QVE1f4bBIQGQOPRlaKceuE59d2PI1UhbA1KwP1OxAko900FrWghs7H
0DzaDum48w45v1oSirdBIhJRBCJ7b2QHDsp8+H6Bxpi3KbgMkiw8WR7KLRFKJiGN
MGcidffuiHV3w6R+eA6lbQXuOQUBIieBIzYJtzK1f3HsISUIL3aaKwVRg+vCsqkN
Dqg98AypE+0F+7fQBHs92/trlDIHnf0ifZ8kZizgjTOvskM6f/G4McppvFRIxUC6
0YH1sOKga4uqlVp1Xt3j/CAoUHg3l1s1027d1sz2sQrOFGolnqe/cAcRyT8tQ99J
vXWSYPYUGK55RpHwes7Un8gBrvW8wkX0BoT/EBr4k8qQ1hD8OafMvatuKUl4vZFE
/NdJIF2BtUgVFFSqWV5zSLLk3vlCpkf+ACok2Yal5xzUkHEEMI+IUFtrLeZIMonf
iH3hyLYsWYmtpA1grEhdoxM8tAJgEyv+T8PYWDzXGHk7twWR3a2amWSdu/6JQ+4c
xwGUK0zdVOjH4wnb5OgBv9wPC37bqO9QWdKnGcmH1rkqfw8Cuw68z2NeuN6MQlFa
5/Cstbxx/Q2tsgxtTw83jmr8bZ/X/IPEgr22gf43KantA++rKR7XMJkUYQh0ZnJD
VXk9pfKVwkNVdtFLjXIYyDDjYP3hF01wvbh8O8hRhrKl1kZhqf0VKxHbMbgm2iUM
7dKe1E1BzAGmJ5JaCNmVHC8ZeGpCr9vuLIHeOEaC9Fs+YpXUncSIaa+f9/95MlGz
aAXvY7ZMtTiiFFsW8h8g68UkpcraSDqh8zu2CtaexK+gYDnbLuB6GtRV+ioAotUW
UaJu4ZfmqXa9Ig4fxj9eS8AtjMe51mXiQBEh1kG0N+613HaFEtEoywbM8cYprNuP
mONClRCbnU589icXGv8DFfgDvVIkrryuQQFgsvhBGG4/++jciI/hAG3JTHzAKkAh
hHlU1NQw82ZN9aZI8E/Q9atR9NRdkJ9EOwZF1QJE0eR7XKsichOJz0juSMUi9TNi
xw9vkAgsa4v/DXMEjaNxr2JYHj3DNb5r5vapOhDki3L5McajbHiIpquMctvbNqmn
A7fRNaLW/1AtUJn3EqNi37O5zbl8ToG+AqkxoN02vfnh18CqxARsCTJsIV7vxKZ+
1GS96ME1aZXbjtNkBdT3tpEtlTpLFWFjyDKrJxB2ietMx4C6ZqL14Axo8JEutOck
S6Qaece8pC2J0M/ja6JZBF9fxz21CRSPitktnJcKRWMfQZGatp9ccVhUnL6dtE1Z
TRmugTlSnBH4gsU/28pHLDt2QhCU03LZBH3jzFwhkkY/5yW1PFUjGcpTHhCAbQJf
GwsFlo5vDfOINM5ceylG2pyzoK6yhvxY2RCSU5t8J/at2+PYjW5/aygUo1oAXS5B
qVSFcpG96bPFNgJcbUgg7teHKkm8FIKdhgAp5EPFF9Qh0ZKXqMpH4eNGgTVmEoA6
CnOS7jgycVqP6ZuwlkWjjVZ8u+BMzJkEj8JO+rcRqwEP7VIhvrRj27pvDTBIRiLk
Mj7Be1LLXj6yP2xs6AiTwF8T6VVuoLvm5Tho2U/wMJrUV/tBdVi7WklqAh5Q+k3o
lz5tPo5OgU/PyFd4xrJ1dC8MlW4DdAow0gntbr3nX/0Zzd04zGTITyftjY0ZdR9H
6EFBV9tUCLHZYZLpQaw5qEACrYCzzj+ZtehyZTQPS/bAbi36ls4cLbj9hrXLEJiF
6a4/73QOQpYenpQq1UV6AUjkx+A2uMqoO7OaFX/pAQrXGb6xlpYpepmazNubLnqV
a3wuAEfSuBjQK40ceoJysxPWwn/4DEh/lvxhx86mIV9tjuAlyy5QL6Pq2eoaS4+J
VGqOmXAYI9AFah20zw7CbBsUAyh+k1xKYeeB2+Yp18MFjpSxcj0zWgYR55yVaeTO
bXeblsVwe/lCPu7B0xZpvxiA7ItimtpX2uaiUvGqPeIiGQAEispjEgMTX35yb1K4
3SFPrc9qQFHP09ezIMCOZwLt6M4uTl3VfbPNy1DQYB85QFYSyYZqWfJbPsSza/8O
iRCqcI6aCxrg1G2V9C+EpCjpQ7hbr3ehmIrjf9Q3EEKRuSW+CUwYYnJHiAsd2k16
nMhi9TaPCgergoFqHfvJcABmafb0uqWyBwFXoJFAfEUUe8ITXdeAeHs8eDM3mrdf
zW4FAbEjGTT/K2s7UHZOvQhwUopkRy1s+rnmj3kHP3ThBpz6nx/zJm1SuMJJDh9R
ndIjE/8hvoObTDugkYoKEZ3T4bVMMLJone91Gf8fwVwpAWGFE3zZPX9EsOiL20JR
SSTaCzfpRU8XLVY9P9GIM9AOqk3xMksfPuufByj3QAUIJ91HIjQF01CwHXIeR5YN
a4g9rA+knsbARYLbufbOON02elzeuQ5Fi2ngEhqJ/jwmzi9bQfB7qJ9timuHIFqD
3QRn4NLOpLjASpQfLK2wFcmIYWlGJYgBlfGA/5fYMIOFO4tfIeUEGFyoRt0Auhn5
nRk+aj/p5Cw2y0Exect8bE0Nu/7+jn+OqBlYHw+OO3hOjWEQF9SGKU9tEdGlqTHA
wn8M6VQzR0sBGuJ8wGgREZZw2uGyfHM7y50tuF7OMiXjikHTtEIu/I93m50V20//
SFq+Qe78ToM3s1KmrPRvw/o5dgTjDDutTVsWiVRIYpP6dFgV0vmvY4FM3nN+Qzoc
sq6MSF4d9e6lMTYH1BxRQBedbcwX6yHGJ5pG4l5ViNySyNQYLRl9yAomeVkDLAzi
8tJan7rUo2dCNIH0zHUqzeiDMCLTXIgpyHPAeYfp6xkSdKmAYyeK8kTIzgirZKJ1
xCpK07iNJCrqfRRRG3G9EqHWwPTAOQE3kgqUuHqJ9SpRuClTnkJphObx1BLSFFrS
4OqBbIVi6Oap0+e6GCztJxz/fORFjq4/w9QqpF9zostVSzPVyvWdIIUjx+jT5Uit
mOjQ+/duimgGv8hEckPkpN2KR0YUsUyGQU6bXbEN3uZpxggudX6EZoEQ+C4rC9ta
cAluh6L3yNO71iByrt+TYry/6f+2lq9Xp3vMamtW/dTmIo+qGHvUIV5BPsBj6yS1
nbpyohKDNt1GknLb5pkNWRoY1SE7PnSj0wGMYS69okKdrvKqwdLmckyeP2+0dFmI
MWa5gAiNF7x17w7rWmpvOgyOSETuWMEL2IlTBMOvR6qyo3OV70o5xCgIuuWywrOb
D04Jji3E/Jjo1t7LAL7AHTv9XlW+cduPKxmkO/gkCVwszbHlACZdEIdaZJBI0VVd
oDU/vpJLqUoLsMm+NXL7gUUBrR1m6ueTXtm4cmbvV4+YU4QGfUpUuqSj4aOCIGIh
gd7TbPZSL5e7qT87mQynjlAtggrTJWJ2q1+A2z3ddbL+1QsYDw0d3gWXopnSz5NV
r+4ZdmYsCWNlpAv4H6KdAtHtdZ1h8P5LqjVtwbd13yxrOsvJ/zB+kBKYqXhhQ/xG
0yrvzRfiawD7scZh+VXo4r0vZvGrDfNzyNtf39M6DCITIFKi0jXlWZr1a/D8YiiD
NbTLgaCiLL3Bw686/VMlVEc2F5tMAq32XgLARuW8ry35OSG3biN9h7t2y0eQvRxF
bQG5j5qow4pQdZlT3PoN678FXK1pOzdlFUx7PfPcOWtjQx7Fm5SV5cTl8s9p3tln
qg/J3PyH/QP/ollCmJ72RFqOt3dTE3gi2nBnuTzdFEUOlzM0Ort2sa3+RoDYUPyv
v33tgH0qbJhH+cg6szehDwG3eysZH0SJhgVm1yEJHUjJxIY0IuPDyMERyXn1xDrJ
3g9kubtOVMhcWxceAT01ptIVOfL+L2rPGRDBstuol8AFkcaF+qhQq8kO1t/wlx79
PXEOtDUbh7Y/oyZSJR2sgbl/Obge1UjmH10kp5Y9TXxWV+cA/mP8/8uiGjyV6Bef
+N0NYhu3/w1PALHBlucrwKxKNZyKHRQTebM636lOPaIHCysNGR8iOhIto8P7xOmt
Tkna95met7sxq2LjOy3NVjxZxnMk5qWPMi68mTV0FTJ95ULHcM40RPgz8wfhO87J
KL2Pn66LIg9UQ0jVoMtLi/t6OfhGgkqUAkV5cs97PBrV166dnXUJsSW3EZGgOmW9
3maa7B/LFBVzOFVqXtdwzj+0qR6C45lHM/0oiTf7mItbX40+jLA0QPvzD+esKpy1
XERp8P3qxLPEYjJFlGWqEgfUOCYeePQ741jL0nlTwVKAhlvuiDXmXvkHK0/zSdg0
Sg8yO66yX3NmmMGk/UbB1ytSautJpXYPLd7NgpjHl/lg2YGQanUeoM14E2paw9UB
BfXUKqMUQZz9Y9kVhjNCs3sb5EZNZx+1iwF+MpDD/ZeKRQGiG7PsL4v/wdiFzisp
HGWzyjc74/RLkWQVl5mvns8E5O59rz60mf2vxMNM82ykATDkEocbPK/GOkkbEeH4
5r7XYY2h59tFZ8QWoV0q/2EnnIX+Kqs1OncOuIv3llX4h3CVcg07S9zcQDP6bK+N
omAlHqzaRPF6uXbEg2sRmPBbnz3vcAihJVsl1MxF3e3VHJgVw/ue9jw9jUewGAEu
gEOedQt2CjpKzwUhYwGZA/nTRSAIGz10McLuVYZrcMTNh4kCnhWHCBGaf862deaB
YAvhJb1x1ej/ZYSVnGNQLIt8wLvamVqEN643h1pQdmJkFOKzUHOyzEUQEyRNG0pa
Jwk+/Btnl880upYjeabCxEKTIUdrTdpJ6Ocwmw6bjID0JxBdrXlFHuKmCfa18mXM
rCB7p7ImYxnYsMxktWa77xVHLx4xZ/xk0IIdegiSXsBEBjD2sGaqSQxOjCmvqvC0
OjUuv5wkc5TUcdedGYS5f0XCAy3OaZdo1U6Qw3Kz+Kamy7ISUe4VZJDUq2i12i5F
JtdkMmE4UM0eYbw1MaSF9nZIsIVDdTgTxcLer087PhDABLNVPtR/OzUTz5/G1gg2
rCvH+AhXc+d3IgXPb2UYV5G3bKCqEUttwG14qTflS39OHyDD/f6UGAPfc4c5lPRP
4CEGO1+q2xyt9zHI9eKnDkuaRrP/s+vZUX1T8BBedemKrAB5OUIUrV0hBHhNxPVd
Cr813MvA46v9f49F7OdfFiXa+DMMRy7ZmQ3dVXI4rpwNk6B6gxI4Rhh+v+ejAi7X
2UuX39kvJkjzioAhkK8d+xEnWoEaX3jBvYQ0UCx8k3Vd6iSvCWfMSM2PRQuSQkR+
Jk6fk11C9/95bJGMIeqjlsO+s9cucuOIhns/UFUKKHMuvOzKbr6DSrxYkZYIYDeU
8LDHqnP4vkkjtY2bHUr+lycRhmJVT93czG2ryR+2h3IuhYZK13s50rs9pgJeNC3k
aFVXw67zlH8+yrYYpsCUgL7rDV1QcdGRTfWLwUBb82+Eoc1x6Iu8autUlujJegLM
G82mjgVx0B/jcOa53OOD+z9RpPxWFM7URD4vyBdbDDt47RZG4NkPJ++j55xVudyn
VwBS7bqPw9Cxq6/N+716cGfGZRwy/LGIz8a/1tCvo0AQOgKKKXZ+Wcm6y9N/DKkX
K6HqSXdtTrGwkH+plYknqTQe30zrj5j698XxIsYYm0IwL0KBPFeoSDKBhFg6HGSJ
y23ki66yRcv7W/BhngltvIMcG5WdpC0P1qgJEvQ+9R4DZsHOoMGb7kO4KLHx1jy+
6HJ84UqO2+1wtic1E0eJc+6Wjv1UlzPa1W2PV6EdqgIiXkXruNLl4tyN/s/BMMa/
MvhCWDc29VxiDdx+vX2avZekoaf0v/D9s1PV27zgB1m1ibIvlsUsaGNQ2ayxiqtF
YcTY1eUBACHli/I1G2dZVBb+1YCEzyXdXGPPYtDpsvqDzbyGfgFoFJnc86+VB5m+
UfTmCs0Mh9fPwTl9zj6Zta4cgzc4c3QpxgWhMmd33wMRdOjen87+C2SBzi1I8noX
ecz5BTKOy+GRTPRAFiV0PgZq2FyQB/FtYzeS9+D/iHCx5ROJLWSoj6YhlC0oU/tD
lNAzPMtktCG0SoRdcWhGaE9vYHYPvC6qU+uU6pg9lUAkzKdi8Da6OKeHtsCaa970
oYouUKU/M+fwrrEQm287vylstIDPjS6BByjYylVpb+1Q9KnAW9X+B80zHpB0jYsS
lfWQdCpfS3+P51VaZ9FdF6mBdtEvUpvKktujIKwhSVHcpTAGA1I/vY94kgULCQ88
DOkCZfN+3BrusqVAQl44OdeRRRJ7ZquhuxujyEajGrNGvbQTszXXQocW9BjjheRj
0g9HAeLck/QCxoQUX1PMuNc2sAD1d/gGhrZ/pPBS9Lbwuquh5IRL1gHSuo5R/z+K
SGSzh8F3WYeC25THjBNb1HdU6eabTMO3otB6MOllCH7PU5iNmUuIhz1xs51t9x3y
YKNTzQwvC1Qvn735g+E0Hb/6D4r74GHkPiFNIMEjzZ7YaXBL+bs49WY6QW+54GXH
rSKMkHllRyN90Gyope3dOxKpev6SOLDEnmBIEq69b/Nb9zSLp4l/MkclBf8zRaOx
3ieMjMgLBdI8EQgUrSntshX8tSNGdTbxw1vF5yem166gbc3WZjmnpOflpUh30e+u
qypZEyg4a2++XI7YYNyyYs5EpRpKCZ1xiDmHLo4qje8vefcN+zGwBj2j5kA7GRKE
eyjifIlCL2Tr2et9FUuS9Zh7BMDgS6y3ABxjTYsJ1gtQTiLUbPiszwv2jvRKazV/
AjHPBvoHRPXlQ1nNRUdj0b2ksymutxU1pB8cLJCyM8g243sR8udHZpb3SawEqXAu
VAXGoCtKtplfQD6eNd+8+k8c1HW5cXOVveIfK7rPtla/c6Fi5fN0+UtFPwDylzyh
uFGfqoKTHhzYZyXTDBK1eiRcL+fkN3+lZqyuTJNJQfgDMCukm/0btwJwNj5i11yh
M6Z4urBWm6gawJY+BcVFrfC4EdTbYR0TqufjX8K5C5LmskAMlR+8DfzE6id8XXNX
iENstI0SnpxGWoCOn5eqRFUhUkBVfjLiY2RWjNjgnvzleq9kXWKPFKZxkM1Q0BQL
mI6rHfk4TzxB2LW/SafsGpy9eOiy0SlTH1nVuLfNkCX6A2jqPQqMxGWd3kpNWewW
+QkBPfjA8gcGSE22U+VXTqNuxlryz5J57jKdgydqoDZGnAAuVdIsy678YnHJrR5F
K8L3YhUBbiSRQ2mJNevjOG0HeJWPGXvsLVg56oyT/HjDYA5Bgoj8vNsRmUXJlLEu
A8qB9JbP7BE/pOmq8GC0853566KXs/cnf6+Afk0r0arpKtQN+G+Zjz++yCOqMlRm
5tf3jyMZu+z1JKrRc1K6K8TF5AfWICy0KhM/K8VJISNNyGDu+Xh+J0JA+kblGMQv
BwjXNDtIlXzM6pXTSmX7JnOIcy+Qe23aKEBNVLaGXiB1nHEee6TcHbykA+cNkgk1
eyJlvhFGAsM37BOx9Dr4NGjpB6Wlmnjl6KTD/qQxZPJpWs6HKkgtmy5rCuHpGXwu
Iwc87iOD5XjB8e2urnh0cRf80muVD8QpsKvFSnX+nLc2F202PKeGfURQhfKuywNa
iTFrmDTtAJZNIrZ29W3onH13y9QYNymkl32bMXHflL/RwoT8BQ5njGF7jf5fIobs
bP4gTDl522uz3E9osRR/WQsFcI7nZYDM3J+pnLtPvLl3/hXdU47z3cQ31xgTuHfH
1sTsdzJMioGI903305doEui3Ckzg5fJ2GpOA7vMCyDcK+u9rp0Lpe1FFTpcrsYa6
bDy5W2sH8glbp6H02HgNTSN5/yhDhWesCEgE37sQ0xkohEjAEtPqTIHXajM1/YFZ
x7EKzuwYDnLeTyDau6CPaVhYA/KMJYCfghapaex1pYxO5jGg1wHDtMvkUcPFdIoM
xwGBO8BNVXD0cdxJavZse+L0QUFD+ef0rltpcUJUR67F+jgyBHnigu5CaBQIf3Oa
mamhfM74PlwiLXgZYdpel40p8Hl4BQmxShL75i9rIPJZ7O5j1PoMkJfu+onCmzhw
IiRNwIs/h2YMLmX0Kjyq3r/Uwa7TRM3g13fH1Hp2+n2jvS/mQwxhXZtbQ9O/9fRB
/aRu2lt8xkqn0Nb40AivdZBxmCougmkP9u2e9549fC5JyJtyCrTJmwu8xKYA6CTr
3WOCK+nmkXhIff84+PfxoC8VBrYUWhSi9TvKkeVZZQJTnL2go1PrOZpL/F9qRc+d
fO7F6hmWbU6vh3wLlrMe+1DWNKgMptIfLBcqLv+nrlIvBXGb1jwocR7ZvLML/o6m
XwyDzUjAWFmO/3PyZC2UyM/kENRlz+R4aZ3MzTxnKM4klMvkZRYtAcSpO5jurl2i
ZOxgrp56HXlkkwM/HXF0pSyYRokg6zpYC76unbp73sJFg9BGtaLH6nkycfqDkD4O
/bQKxvDlp9718I+oipCDDvToOY1OwgR3i13Zb9eqq0f1W9kOhLb+9McfUliEseT8
xnL5Glb7TWt6vlzBh2rco1XC8jjPQGO6R0bjKOxD0RyA3C5N0aEylWbeMugZH9is
oKJRPBzXnlrOqXedEAhqBBRD9qG9rvT/u8grO9uUiaJSVNIAj1eholtXBnByQERy
HzjiEX545g6d3jOYNefsqpi3oUpjVdGFT143nXzbhOU8b/SNT9+HJ9p1lOc18V78
ZQWNBihG2r0TId4F798SeAbaoGT7EJmwz5rU8aR2IwHi040gCuwfasKQWH51ZTIQ
+mAesHPC09tX+nl6GL9k1zYeK9dsavSq+zYgNpB+/aVBoVzejMVy8rln6ixsOJ04
bOXc/4S4uuGzD3H+Z9CvnWM0JewO3pAXkUXVNqECDaXi1A2k8PREWzI1aq8Niw1x
P+eICVspmwVI34Vy49tBzopgc+bpB7pBzPmXiPMiTnR9z2sNax0ImxCa1pVdHA3v
QMr5HHPuYcxO9ThV6dNPFkPGEmZJtDIhoSAuHM1z2Pz3yGCiuZkcL9k0O9tkfMv9
NvWkW0ZpVVa1er3WndDYtpw3oAMRJK/lz/wXqCmYOXHxB4h0raVGDIC/VVRnKhia
xQ1FjtNWkRLI2fW81xC1mWb/pazZ1tEFpR1iOF+HRsjR+Jix+R2E4wBnDF8xdHUV
UsxzlTbAw8pUY6kAH1whVHSfWgQXhE4unzFGUVO6HrN0P/DFn5Faus3NjhhUuRnd
nNmPvrf8jUH7hmt1lUErU51b+gVhijBYm9sMVnkpGAM4zcZPqSO80H900xtVlL6z
znGOR94Gn18nFK4rpzXSFYBdfkNjAUjQKhg3o2bjY01tJ94fyPIa+eBE8o3oOK9x
dK22pKyL08ZtK5Is0Jnok5kUGeBHk93+NzU9DyMkCt1hbpha/OCoGKs7l9ScVQwy
bu0IFxVbOStc8Q5ddCoedgxiUK/kwc95pLWBUJnui1Y+Dhl7NgtxI3jGImWdC9FY
Yu967BEAFNkBHNZExFvkZEbPj129l7/scZnVPxiZ6EYSfnNPI/60pAd7I2tH6rjf
vT216L+uEi8g7D+dPFKfnrXI/FntlrB+Jr2Fw5hkizjP+N38C5DX5dx7D4DG/57C
wVcZcplQo7sPhdWkqMpNHDH8njqRCqBQFdU8ZOF403XqePgvNIinchUSZKf8RZ7B
gRa8BdHbf2j7zdYuMMHD3jmg66NXbAascfHKG07SGRPGUnevS5kqfaV3IXZ7y/su
lvP5PUodU6couEJo/LjoQ53YSstSpSI6//304+ryVWqLkZC/e6so7w0YIWBUsFWE
VW2PtqXST+XVHkvUa1NWAL6WfaWWdIib49m85x5L3njd9Bs7V+1Q4E/lcrUjykhb
hhQrj0m7rbwNRu37m9RRlW1gBsF2SbNh0UJ86cCvjML3fOXFTPHp40z60/H0bbx/
Mrpf1Rymq3+hF3lYAE981/mr2nHpofbNbhckdybUeiol/ZMjyJymA8vTxaYn+oAC
Q+SxMD4ByHqyu6w1mOXudwUX1CcDBbjpU/YtjTpzftRPk3BxXdBeffQW1dZ2qmdS
MSU5hXc8lNi2jymckQTrLxh4iIfvKtO7B03jy3W2MR9jKR+BMV9Q4NJyokLYzvH7
W2GfE8k4Clf2QTCTHQ6ythEVh58ASRWTOJi/mPae09Dve1RgsWMd6h0cIPYVT0Kp
wcBVonbW5I2KzuYQorCLNGFvtbjcy4/FlTBbsjqyjoXxNJdcGXyNhQkxgKq5PHMC
FMeARP1Pi01sKlc/gA+n+6GxBtItnfEPJO+AtJ/Lw1gumCJ/fKizY5vJzEuajyhQ
uRIymaYW202XZ5fJk6o2jrbJR9+BDI2pHEXgL1sGlvM7dtGIbPizM1+V0RopAPeU
5nNLPO23Qj708DvWRABCVnMQ0hqrUFK71DHBAvObwMLqBmFUFUv80lXda7FI8/wt
Alx25imUpeaZHyoEP9gBy6bExyqHl/2vBLQxdSXrtOOV+HFUIhX6KxT0PZvNcPCU
nM2lh+phOI3cSMVosyfZRNi3DDtpkHXwPDIOVtuf+PkMJ41v4bNy9J2nLIMCwwCT
W1Z/KsnVUP2Wy9DyZyA3N0FLyo4pQJlfry1wboC8nIfXXsLDOgL+Ro/1ozuzOSXy
FuVKyNzgDND9eW2ccd2LffN6Fmm/RWIAPnKqeeEIqGTLKxa4zeMBI7bd7f0VVizr
/+fzkzE8UAds/XaOv1vCfEUWsb7Mr/4PfjF9JsGZaEQpSEonBOsTlMsnRCQBAwTb
Obrx+kOcmHJZIbKN6pJklPZHErP45ScLXJIUGZkrFo4/GNe6uH9Vo8NrS/d2em8z
Rt+DMG+OSjuLoW4EX658Jxs7yXrxa1HQQLxoZxdmTuBDxsI7l/vImLD1s8o2itO7
03xZQ1zs9rOmbYBZoc/LO7Er6wST4X06koslHKjCJifihnvFpjUHv9iQ5PsPatV2
CwnLD7SkV2J8K4JcAqImLjblhbf+jlRHoujyFYTRfOgEA061jEDIi616K1Gg14Lh
P8fvBtdrcMGcD80cG65mGjXlk/6vzcRDxvf7CFt9Wyb5tzlFcl+Z+y6w3W1g0cac
pR6SgQut35Na7x7lsfuzsVuCzCiAFxKcSBTUt1gikczOKPqWl8D5Q4o7MdUC5/6m
Er5ySYHVa8WZ/Vgyef7R/UjtQT9U9VKXfUqGgmgGSoJw+A/j3NPZeyyrYNHF6Yf0
7ws2OJfTqz5OvdTMRf/Jao2AyTYNaPs1zwoaciMqF/nkGUTMI7E5XKJJsu/xK0Ps
H+Dbo3G8Spswki1LEOGPuial7FvVGJtIUkQTLxPX89aSViP3A1ztQZMVCkt3KG1O
t2lhrdtrY/16zqqliaI5AI8vWSQfL6cIRnchwGaYTDmfpO5XUo/JP5icOfndkZBq
24tp7I6DabUkIvYlzXW/HrQPofUbvS+jhBwMhX8j+L3nxK1fMU+TlYCUKE6gqDg0
//y18ZNp7gNQRim3NYW3zjE8H7fQsAAAJk31wj3MNpZ348yT9C1HSy3c2Ra575Dt
N4TFymqGx675R/DHvGmJ0Huljdnwvi15khd8v5Nrj4Vg6Ij00laP+48Bg3YTf4vQ
3CUqB4JZItykWey0yHDrrGRfPCdcJFBeLsvt+qZQ7EugWCSDABu9tXqmSHw/gqGC
sPvNfOROKL2176au5JT4pMa/hjU9gQJjMdtq4nHkDcpnE5VCS+//nt5jwJV9yuS9
bmRRQFp7CPII1grRmj5p0IOrVEETjGdKpYJ77NqORmlM3FrUdS/eUK1j4Dz91rwE
xBcL6fiQvZdEr3WVEBfw59alZhw5oDcSm6RlQjW3awVxZly2ENilg6KOP0y/HtWs
XyapDvWXIoCUGqutIaGLtH6ljfg7NFEae0zs6dmc8Z944X26hm/3vQHd0aj56RCw
vwcrljQxohLg2flvusWdpj/qQFINh03iwwJVDwZn2Rzw8v+yhaBUEkPMpsavrAsR
PVY/8nUBfF35hwjNovco4yWSeCjkoOKhNTVD/QOkACq24BIPTHYz/wVK/A/wFCXq
LKOCu24ix4M/bJeMKs0/uN6LTOsQWBAXp6eucIIQBRD4Q4QgyIRbBy2hvytY+a/8
yMFeSoQMoqOKKDyuQh8y3FzYiYY+sdFbcaGH2g6cYyvaJMMAyuu8zle4qKFg9K3A
vz0qHNzwjXdvgx25pPh7DRphqSIh+kDi3xnl+rQ3s5oPjSM6cmREDG0+BUhDYAX0
npiDi+IlJganUpHNA/EFI+8SUzdQlqVLZizjZ5evcG8G5ajNH6XghB6p6uyaO1fT
GjZ9atZSiHV+fV6A7uBPfSTfLn6J4Hohwotr0rOSIpCTBB0SRx15zq842pVzy0Wf
wX6/ASssRtAh2NPD/H6R7y2T4Rf46afzS/3nYAmYV1y7M4vn8pJhv4kHBChv48XY
GsBunIXcz4PyOrzXbQdzK9wpz+8LqgIX4PhE+lcQDqOv+qB0I+ql636I0aA8VOD4
IKORjlOhYrvAGUcHzKzLukI1EumW53Eco8pvezT65qLcOXYCT+WWyeWQBQltukb9
w7deX+UmNZiWu2WifX18L/g/4YzBsrnzZkwh/OKr5MBifWjXp5ZgHdubKa3VkfVt
CkxrsjDJKxFqeFd9oSywWQAG5GEwZiuFX5zck8cvr5BBJkks64o7n38Q8JczSNe/
sK3IP78OjERF7781cf3pUAkuGljhfH6HY24RCUUa6IsSYvh55/8GcSP7TE4wS2GU
l2Rcq49uWgbRhBBNXTUpfDcysfcBSpScbVz9xQxSQiGYrwGRNBQnrBNG04rqI5va
oYLehU4v4eYZwl7Obgt+4O6F/8UlWcRbc8rs/kgQsraG0C6i63Kz8XeuyYflzk2N
UiT4NvwdC8Dl/AThyCj2DkHS1nYnJ/ajlNbGg73Y0z99ywREc/yl6uZUrLyBgqs+
oQawr/9deve99iqu3we4AzHSPITcuMJkuoX9ohuoZGlTlfJSPAzrV6RHDM5h76jd
qdzMAIBydfrLL7BkB+z7MN1uB18lAPmOWHVuUeAcLeQzM6KPbH+kYLwFNBv0aU9b
mlDuhHgXlYe77QIW1aCOyKXkEQnzLsR3MU57edNB1DE+f/L8FBEZYZihKLhiOolH
5Ol4zMZZ5yqo09Jn2C+Ez91mEKgDTxmMG+Pct5v+OJMKA1Hrzs202QIxnTDBeioZ
H7nBZgg7P0Wm9rAHSwfNiXN8NGg4DZNB6NvaHsMmujsJzYmkzxTFeBJGCsmnJgsu
J7Osg0iRhQEQUNnecrR77NIM/KPnsuOQA9yRp5/xW40RzPhYtLtu965VmAZevTB/
ukeO2bsY9DmVGnJaoXgK0KqUhdLXyKaM1tIwGGIJrICjuGUc8IYakoBindybM99v
D0aLZdzwrRRMzbAAOwGmo7OChtoU5mQStsbHk4DI31exdkwYdSegdYP7Kn8Ks0kB
lMkFYJO8kW8qJ7TIbOgBe2ZMLKodGsu7+RuLA5itCDWIJ//m3YYfaG90G+g9nxLR
S12vqLrzCASRTc4CjrZllav+7yKinmmBNMjmrrltfviesqr2mET+u3EnirVql7bI
XqjGOWJ3lidgFErnR5YwnDAPy+cm1RlddrKDSDKVAtFr76LmY752ue4uhYFNOUCB
lDvjRkrSma3k0ccaEMSlAbQJtPuLqk4XQHGzhcFbVv6SEJNVRcjE0d8MV1gtAKlP
koz0W5Gz1cfkAaxUjIlWVksD7dlzX+JBQwz7mo364b2OcQzKz++1qytgTNQnJMmh
+R6oypeMy3jDPI734xYtRmUcSo52T8jNrzSh/V9LoAjUeDw2/EuWSD8ms/eQbbJ9
Q1Z+skvW+v6axvdYUSzf5GkdW/sj74tNkYHiVMWZMHK3HwiYZ+7BFQkbOWy+m3v7
a6smUK2RFMGuoZXH8JuJ79IWYhZnsKVR7c5GLt5wcTSbd/8JRorzVgewBX0H8reF
3RmcyP0TH3XUrmfPW1kUGTMVkzeIyYCDe3b7qQEWj42XPo+o8nkWHrkHtvs3MllC
HblSiibNzKBbVlEYfODCUQpp4RuVyL7Pg0+Esf1Pls7RnXi1vEh5j8IuIIMniDUZ
+rnPCzpPZqt1gy7tSNxChwDTMXNwQI5qH103Kp5dEMO9s7PJgV0MomTObkAHbTCl
rnvd8lhjQbjv4HT1Dv0a1H8ufZAQImD3W6AYwJb2rtur4kd8Ti6NT+0jYmEcGmuZ
+EvuJ+N6dwjDIe9Devpwr/jPSJixyR7OR8UXdX9lCwzkTyCoRulSP/dKLWk6wzeK
WTimxKGSmy4KaipHqQtOq3Jvbl8a6aPX9earLCtEhyAaJLKxm4GU+FjK7KYc/8df
Kx6JeqSw3zwVYGyklFf3RM2+jrQ8Dcip1xfhKmvFMO+4dnG8WR9BDE+QMQIUpBgt
DZVdpHiyRGm74ZGoKk9bY5/NLxh2P4tJpYCs6+OFgAttHoFe9xlZY8U5lHxbff4U
XINvvdGgP2xZ6GYYHyxEbXgNav+49+MxGqcw0F8bZSNVv4zobHG00TCEBPRfsz+r
Y9kuFQKc6CBojZ4DvVvqyyVhEKvsigWk6z+cOt2qVdlIUQBhV/mEsnc2sYTlKuiK
MaKqH1O/nTeNazG9lZrQTZ7Xf7Ba1KpCfSJ1wf3EILmgeKxuFKWTOFBqbU3zjaCN
ORXHyQLCnjZ7/Ndu33iceCIzRG2heImiNvhiW+mfPzvxmI1t+s9utIwF3SLmwLjm
1qJHXcfox1x/yQW1zOvIa1POf/xwHccd99bPXMuAR9PhcN7k6na4DK2mpopxHIga
+MFlxU9gK79Oe2my7gu/KAD3zGlM9tjzMJF6QO3ptaysuZhUXnkKxY2xEuiepZCy
hgFba2ZYh4nB/7f9foqJ1n+PRIu5ivGta3jaf72zEx6zOv/CDJRjjzD1RhrdF0vv
rTTnqNvynPJQPGPbfDDzgYmzlNEnkP4mzm1RoDS8KqZDlKj2K//6q07Z6YN49p8o
38qKGyWydEHXjDuZGOnhvMf0TP1OzUa4Y31l+k0mKEQDlAkh6hQbfA+HYPiI+HDQ
FVd8fqWlo0tvjbImiXDNDY5zSzXtzeLlOZsP0UfAVKCXkKc5AjStfivTaEjiuSpO
ZDiRxPBxI6oCUDEl3SFI+ZmBhOECH2IhTo5nLnSGnFXN/ayCiHwRK+J0rKRki2Hh
EvwZAvh2u482V+e5vLoDrVXcgmUqGy6MXWuRMP9cuYB77COh+0xPl3obmE2IqaX8
3doTCA4AqGfB4e4hw8L+wvr1vEOzDzCBLLQFaJhVsUJaafxrLFPaEQYliDcQ6VAS
NReNoryJ3R6mLkbeWyC3N+X/nXb//NmgA54pOZbLHZS8IHUJn3yvY52K19NqbpuA
W77rpWV2ZAiM429a/bxjlB3VS8LddTPsA04PO/uoQ9DoHJep7A3lsfwIR+XO44O2
3d9yqUUIH12gNet2WnYBInbxdWEHXLpyOz26S1LNy9rdGAg14vDmNS9k65MSi5Mx
H99JcTbg+WUfZMcYnfNWhOGFDrQ0Uo+Z2/314nUaVZpIl26igg2wIno4g1KdzMeY
I/WXly0S+M30ruLwBYuZuvek5fweQo9LvIMiPS+++KFO17JDgK1RnAO+uAzTi5bc
eM2y8e3bb9uW9bSi9leERw2ZBIUzy3CGrahPup3JjXTQN0YULXOrNoFLJ1dfsXZn
BX6uro9NN0ktr9CwSUB/rwyDlLD/Pq/TYD9WOHHm65jt8I9E3qnsHlngPQF5SCX6
vkP/9pXj9lZjLu7DSfScnCKo/rypIvcrWspSD9WbtQxRdLgnsZko8pWbjiVvWJbQ
9G+fMZwKPE62sp7sejqpBbCS8XAd/9DgZejcLf4viBogWzNPUx7HKmqYPMX3WfxN
YrwwkkGbNJ30k0Gf6el9RcerGPPmi4On++ovmyhxxaovR0KemNDR05n1xZvBETd6
Rpq6x/eO1QHa6c1gG7JHrkbH/ofbqEmxy+mru5VGJc9f/JUrlhVy21j2Lw3A7Fds
YH6B8+AxQJt4qYmNlXrL/FnFNIMg015CCtKUjFhm7W8ta2QoJ1o15qkQkCAoO8K4
ByXU76jFYDPqAAvXeS1qFlDTWy4VyJJq+BBG0C0zss2zI8jfiPVEHG2eyorNLnSu
x0/Y4nBzWuySpQwpCYOSy9l6DUBHvnilTJ6mMe9meXk1G7yI+HaWt7etaj4GX9XQ
8If9ubo0ssJZLC5dB+12lmkCHG+1le3tHDyMrrY+TJCXoFRcssDLOUwph6GTWtlb
LZyBLwQuaroxFX79kjGL+9aGWf0qL4CKN7JVbvZRw+bGsAJRQJR+CzuPeLsZMdp1
ULKDbApEfjJEkgUfGcevu2G53L9zsIknLMzZfPE10Nm4+oPAlxJsjzJr6iKbOi1Q
thOAn2+lhwm8JaTvlIpcl2QmvlUKh8c3Z2YfLaqyZpJhEgNNAqbS1ABpEDSYlTCC
9bWQ/HCAwtDzRmI0Z6aESDGap0ym9kB8664NZV9QIXlknkWkettBuAdGg1JYMyyV
pXPaUAzKjNfFeHaoavY5MZ78PtB9qmPUEA31xSi9YZz1I3DSDCPZ4TJZhT/J8Fg0
h1CWKgV/pIfS3DAwFCPi30q4ZEqMW8jnrCj7ShklRE8S40FRAUNsVzPh/CLxBPc3
UXfwBr6mBchn6JH2AhIyqeItw3O67Ita96accI+e5phffE/IsOyxsGFOUnCptIzw
n1970Eq/Ul0sEee4UYT081FCk4CRyH0XFaHGpqFYdeptEHrTzOTno/+KwolS1RLF
Jcc7GacZa9yRKCLPCCIERGFWgHO7A7XW/OEXTX8AB/lzkj0tB/DPFJ8WL4ltAlOK
inMplGs+ji/nwZeejX6ZQR3aSl2VmM5tNH1OI88wdj9LB5nEplavUf6dgrLaeDo2
BECBz1UCiHqiFxHXHNHz5ioyRpORlYXFdrDkHS68kUOodoytdkybePMiIctyghk+
r7/Ww9vQJQ+PDgrC2bkI9h8BBkcfPJqls3eoq/82p+mc8t0+3dPH32WqaI9HbG3G
+mPwEsFlvy+OQq2EBqnwD9wS3bINVl7uCHVMByzVKvMsJB8F0qJWIgRPqAS2LGRT
9kX8vgzIwMMFhijt8ulMMKBNo5NyY7RC+HjSt6sbnSH3CdhztcRToEPqCdUs5Lb9
f4b3V1jJDK6WlOHvz5iDzdnGbb4VSKTR/ViKO3bmMzrt4TtDNUDtkE3Zj513o9if
PRP8T0zQhZPoxAeU7iiF1BbOOWxzzvTFU65QrRj07GbkbBgGvGuLYq23/0qgIqA6
wTkEF8Asd5Cnk8ikSMhp9F7V1H8KtrSUJTGXwvu+r3qgPjHQMutGdRVfG5YArUjm
aux15pdaXg8MPjuJyB55CRsbUdZK6n6yJnsc5IL0AMGn8vkrJr6uK9mmylz1veK1
Oq8kJKPMkkQZPmqAz5Viz/n+gtIegAQH74pT1WKrVEeUry60enr0CK3+UU6TFHdn
oiWYJm3oARx3eQ7aBYV2N4EgFKzjWc2wz7sO69DtGDcavCyVNzmnilx0/bUW+oxu
GnoszAnmUnJcNKPl4luzSeB1cJIeXFrJfcFQ4g8q3r3BdfEPFQ046zyAaaqNeT1F
xz3DkD6RrEMTY20O4i8foOIBDbLfmxAkZ0AfsAbPYiOupKYcoTNsHHkz+0uuAm4F
Bs96cWYbeCithhIrOcm4PE5On/uuEM2/BbbcjEqHsaxp77hPo8mGgyoJmqSxM9Ba
1Zx2TeQdDzbAbYK2ViJAQXkPJ/Rp2iq4abJClcwl97XAOX7f0XUnBF2ZyVcyrLFg
N9m1zUp5KiOKqwmd36xBAUcrP6bG+DUEvf69v68B079TPoTG39GPUAn+QNivVO34
DChbtNcGl7SUwiAyacFsBoDLna0pmiA2m7JccpisaRzw2agatWlyPw0eoPabjSxm
9Z44kNlqpcRRiETiLPlLaSknBZ6zqEvAyIZxP8/w3WN2CqAuwi4MPKhIWwxXI0fa
8QCdttfl7f1g2BO50ysX45MBSj4HaBBFdk1nwZD+oDQFKAmlwLfnfD7mTyLeTW1N
TJ+83rmtDVfDoThfipYqF0oSJOw9iKHSqgZ5UPWC/INRiNqe/Mnc1OhpKI4qdvgO
HI2NtxGxN5GhtqhM6iiJAloSCO6ygdULoYnj7ajqUaY7r9RLc7IibMoNjnXuvCMP
hvn08KMGM5/WEn/J5FEWOt3OKMIFIKMO3dOfQgtqWjAa9+3/krWehn5uIcF5l7yw
TCJr1IzIkn80AOxDng1qWHAuNzXsF1d1qmOG0eMcmsUxDg0C5GkdqtYOLBrdCGfm
+QsrkmBX34PCEqcyTIyrI6lgahz5aTtbgd7wQRUXMm/Y2+q7zURNfEXTNPaB/Sng
AzorhDB7hYQZzRAu7qRQ/6IpHrPtLevnZeaIMgKFa+GGrYv8Whh4Qajf3qwjFOto
LzhtmGGVkmehO+k4luyYn8a21Kv7AbyhthAD1h+8lGYozAS2frl2CSpPPlj+T/Gt
M5dsPK+g0+bG0DEDfHEGIEH+8C4+PZ23d/ULfqYS10pU1Od1kAkc147jg0q8rjty
RUTTxsFwxYHuxDPpRbFMRG7qYhVKo0STUiNtrQvGXrSC7xkxQbmbOpmgXG/4DSdj
AflGgWScMQhFGd/clCM8zHozfynD1JFcryyI6JGEsliv3W4gu3sYYZnXHh+vE3nj
wkLVmtG7MwQ+NqV4FNSwWXBRjcTTHzTkoUEcJw/kAIuUdET/FepRWHAgrI42LAkC
qGaYLl+J/jgbo/4+VqZmjsV5NTrJLEiaYtdJ9ddmUYC2QQMfpcAUUCpsXgTMbByA
+ou1K2/4URUujlJlcVcgyJRxV4qHmnPNDxSaBThkBErGwIjKEllR+P9nKy6DwSaI
I0a+SL0lMvRmiLdjiD4Ek641WLEDJ0Zfz+H95L8xuWZIGzMY1crDp1bAbLFwitkP
WilnjVaw+3e+E9daF9FHhZh9cm9uba/DmEiL/jaoIL9z2Hm+Etz1Xt4Kl0wBN1eO
xVtLKz/juf/SNFFlDkhVyd60Jx0JSRJkOZPuI0756kLmmCVeYsLIdb8bWEc7ZglO
1Yg5y4jBL1hheHCQHF1/hoRrosvDGZS4jLP291Ax0sfELu+VlIdYSWkcsWUJU334
GVnx3Nyz4DDhBxD3m6OgQBWGWvNMuOJzM/Qn1a5M+6CNMopN4yhIs60EANItabr5
XXvdfbBwOvGdBNiuCW/8AHfNPlM6bAObRVhd6+vGXW4zv/ed94Qkkcbq7zNwuTTp
egyLM7raNZB5Q47Xh44B3fjxEaEuQrprWDzBy7kHMvKtSIXO6nPkvSATEHWz+uGP
igpgW6qp+FbjX8iVOvKtV5F2VA5g+fJcpXKhJC3Nq/PAxjtSQcka2KemFM/tcg5O
5mSuYSWZSld6TrNq2bf9LIvZhHeVnfC4MGi/6Dm4LXK0L1con/ax4AFOB30zBN7d
/UKoK/hDYxAnKxXu/qv9q/DURqrd5OGTT1MdariV+XAwPoacrMCN3JZyDZiousGw
1xPhZt6NALBJaYhMGlo31Daz1Y6f8m0tb+5hNpjZSlUrvodEjgROyAG1AHKADHiy
qPJbL0Ck2O+fRFlx2smdFvhvNKhRb6BxFVgh72XoXhnVh0zK1V5Wz/UUGjZERM1l
7g9gxJFajSD8VGY+UMTAtWfmvSO+PvfaeVdAAAkj972PsA0KLmicGdEvJOSgzHXk
rp3VVxLee0yOHPOzDLzpPvhcqZvfghulusAlqSGseLz8vnzOKW5ntRGQ353y2waN
u48DqAX8sK0y+3Eo6fD7XJqhsl1sVFFk9I/9pCsfD/9skSI1PmDEctqqZomeCSwI
CdkHs+BK7IUTgyVUHqTB8jrrT3UL0PWY+iEGCbDgLl2EU53ieye32fX1YSYtPQM8
AZd1ZHtr2aZiv0K1tnBcze2EAwG6UzBtI5g2/A2vVcUL7fudACZ0sFVYZb+vcH4S
EmKlThc09mEFpZMoKHgvC3wbuyV/NMCRYUs8Dh17DutVsoN+Dqgzut4tCWLe7YvD
lMVOPysEPakkvMdBoK04Q9hvn8YXUH6PjtuggeSoqi9bbfuZX9NFB1rvQYg/rA2w
E1GJ+eI+imgElyz6oozxI1tuWs4t+X+J4lf9xh05Uq4RNMLt9xYQnNItuIWq42Oe
p/HTLQk1WWj+UfulXv/kWGf4cl3aPQtngrOgYK7Y9p1UvNwWn29Fy8TMTf10oZSc
vmksamQRXxLyGrZlLUgc+ozsRD9nmrOiSflSod7p4jWlPROPwM9ZmZi0zyDEh+2Z
aIniHDkiqEcm0GeRW9aHXs5Nu0W5vZ7h6DFIrgTV9owGym9kiI2QXGldl6EAbHLI
mF+w7pzUCQFi0rpuZORsIqSBRW1wi4JNVpSPjCpuePB06C/sdFhyjhSOhDj7r0im
I3ccA8HelHJSFnytlFjxWyiU+n9nkEwxgzmD4RsiIMSWBsCSj+CEtJfan2/S+P+p
GL93dh/eZzZVctt8h/NgVOIG4r153bTokl/gQJix2F8VQ7qoqVD31t5e1Mw0ayVH
o/1b7VONIUJNjtirv+eVIV4oJqjqBx4owCvgD8ThReILIxEpIh/GkOCCdHRsnx0c
b7HYs4GWq8BO7Jpt23KcIh5LSh7nNEVSoB27pTUvPybev8Ec+NqDO0W1pO3x4GYK
8yMb8fAKAVBZn08x+jQ3ja9NIGiJWghUArBo2hAukW8FtTRks7TNh8PA1VXuY5NW
+JYN4QKjqOF8O9NiEti/J4T1R0Ja3bO1bZRdpZLDZFtvfk1DOaiexa0LfiE6wGZB
Zvfp6XurvQli1Esk6Q4649VkOsvuwiCQVpqn1fVnJFy4jCdx6BVPNlbVS+W39fi7
xwVy1TO68F1reaspgrZTigAEJJyFHY+ONq2RgPGo5AyzlmpnmrYJUQFw/aG8Po3a
Uq1SrvmQ2InuRydOojZrIpsTMmZbPDzWs1VfS3L+uAj4g+ulPUwW1btY+sXQxq8t
lX6dfsRRLKEC1wCDDJTf5pKSOzp+7nhBoj5x8AumJ+76kmKLs2I+uEPKX9xZCrjK
AT0F7BdnonvIXkrvNafOo1iToj09hwwKIyUIk2NdiXy8zr8rwcF+FocQTtljC9+k
tGq8CzqY0Kl/uPISSyKjDhTxZK/xymJlr4ATI7P0ZylU1fURIf7SL671USLm1Zog
P/w1OwdDTcEMgDr/ggh/tyVUJLAy0RQrZUOfnZKYsQ3h0Rsh/U0hUa0G2LdQa04l
CwigPo92rkRQqT3KVtJm9jUQCJiAbnUH7uVDSQ8rpaUJthAuU6FpIccJc3q+p+l6
BVZigzzKPqzWCvyaRcX3eh5UvxwGLqJ3GcBR2niyo1DQrYDpK/8ygTIYdC/mCTCW
ckdEBgo6wFY9v8RndCffbMAxDyn1uvJzmDheAVetEai4f1W0LHknHVTkYf4w+0h5
Ntf6X1eR57K23ls+rdCub5NFYq2ibAvb7R+GXbZB7UxptSHP12JdTq/0hzj9Dnm3
L+0lOcrQJy3bXAC4Zv3K2rCUJLIxn3RwuderIA4MReWr40jCXflvsUFSC7/hdW/a
arokJiMFVyW+INHU3CbPgrsANfqbUhCkp4AbIAx0FBos2W0AAbDZ8aDWyo6PbaMc
UkwcGQnr7FI6edv6etmszFTP1booggKYCrCIX5YsE4nH/htWH0dOKYFSci31b0jY
7eKYZ3/MYDNsK4QtvjPJDnJmBiVvtUqIleTRX0MZHmU4tfH4yrGnio8BRHkZAueI
w/Q6Q4S/d8p4d+Fmad/eKh89L9JdrfFD4uX1cXfImZ8g+cWLWIA/LULWzD2cTnSL
BLJjXkH4v0T4TS7iWx7PshUXNipPfVQYLYoL4iGeV/CQH/a9JGTmYDda9XLw2yaU
raAtPTRfm/NPZ41Jphs3Ay4+mdubTT0I/eGyeaPpFaY/+eq+TW0gRUFAMTAib7nw
PAiia7aEDFDSj5fOlJJFOJWsE1Z1ze9b2tfhFSn1mCXUi1EWpsEyaqNZNTyYmxrp
18vQydDqdKYrYw1xGyxxRXOWh+gPoedSEPQz1/NXrmY5Y0X1VM0n3fzJsIsyoAEc
nBnRXFEV3qciy1hvlKlqklaPVoK4+1KkvAzKpEVTFRg86hL2PiaC2khTGYYAmhbW
bRpXD6Ukve3SQc2mw8no/f19YWHsU/VnjolR4gI+xRNGVVJL225WCcAErQbxfSyc
mk0Y/Dy8K96Hut7D/Xw/QotYJEyXADv1iN/ddQdFrCcUArJdYRS2VL+M93n1gQ/L
VC1aOsKrZSfYPgv1+Y/hFypjgm3OgKV9LzZJ4PRpCPbTktN4WSEUgvJoMC9Dz+3o
TjBt6wDS3jNnSbNI12pEoREraqCP07taKh7yDTswmkl0kfjKbl37ppRLeOTOIXtm
ACwjTC+4+0aQkWDZ2muPGHon3i3dy2BR5l/VQ8NC1iXO5sXie4tOvsYi8DexUYYj
NGCZejarVn78PdEblo80KaoG8LBCibF8u7zOkYCPzvvaImSLGjj7jx0ezUzi/nxF
8fPo3sQA7qAsbL/U523r71AVTJmjQdB1tIFG1NNgwygv84hO/CbdC/j3mAzupCTE
C6m4OohWPDzHkOjAVgxwYsmH2rd4kMWogoMu+Mfh+x95so8QW+MefxrCpVjEirQR
Bg9mlqLh7xbrEbYfBEgeyfi/+tLcyQI6CvDr1ktwZVojh0//h84RzVUpnXMTS1ra
II9pXP9NZ8mmG6V2ij383sw+lEidghgjbzaTQwZ7ssPhoOA1J4fs0rjaRMpTM+47
SBM+3wOZUERmzG/6sl4IYTlhrogvX56bOrKNFE9pcWAKdMWP7GXFg2864VHOZlb9
etqUl+gL75EGL2mpgflw72pxYnIlwk4FJb3AHbptT7LLJrhW34GeNfDxsSSFtqIR
zTHThOMbqoMM08oUlujK/UNYQ9V2eyvFyvyMJKye5AgKK4F3OczjwCqWh1++k6xH
ciepCRLcjZQigbq8Ykh15T08uZOJnCkhg6xSvdIx/WUi08tN7Q3yR8OoW97oD42h
Jyu5WdpsdI7EQk3qpJyUEqfeN1cIUSamugBY+49rHw+n+Jrg8SqUAdNgAOZFYGea
5L56ihjkm0NpwX/IH7QiVk4kvue46o+NPMM2wK55LnsBA4HKqLe2UnlgzCPnLf4V
2MJxN+XXNj02BggmGIEp+4CgQfPjE7nF16rfjTFCATyoOAXnHL4Ub7eqafr/WLVP
4AlgwFVBxmO4Mm5Fn/QQ1r2faBMd+Bf9SRqVXbBrbtxcUjiC7fCKMFAQjU0rS9Ka
e0P1XtmxE5hqKtnD25iEZG0Tej8mRa+gMj+QhT0qUIyKxlHJ3nb19uRA0fcoMbtE
jJhYjlyoUvmwv3Xp3h7fmN0sIL4e1+4xKEgpxshAqo5UerMwT5Qrw6P/2mkxkGn8
w62OFG/yGm+cqvtOsIYZaN0clvr4e4e4kifNbDilQAWXWZUzuYj+9/eSpfLOlL3A
TNTW5FykyXgwoXA2NhH7zNd/ZwGT2k/drFnZm07wbgtTOTQ4O3oRmOQSUE4YbAn+
SQwnpj4n80BI2lGisSQWtM73HpyH8kPEzcINFHclkpFGpyJh8MeZ3RtdbOtlIaVF
S2gX5ED7mNmsGD88mWlahohm8Rom1QNIW2L/lt12rI0LE0Juj1ahk4LK0SrIzJFE
aYwXxnfUGMGgzDFROwyaVSoTc6z2dHkAjEg7AZC8e/0/2Id3DUQadJ6onujI+PET
/CReFUcdZjYMR3xaRni+6D9VA5kAPmIuudHiRoc1m+JcUHiJ63zvVwsuKrsWD2dm
fmuZ2gOmx9GWCO6D9fPBY56tp9m0dCv7a4iFQc1XmpdJPTWvM3CyCpBGBnXm/+T+
P0AzGTmmlH4kzU534IHU2OYkH99IsKKgm58LavloDXqmoOYVDHD1iENwkbMk/zJP
BKgptaDZ8PgLtA9Wr7teLsTLWipg2GFxvuIdHGc9WHJTTGbpbPz6uv6LYCyHfm8f
vvIYnFPePIUKKakr5l+rkEK1q1NhKNZ6LG2XC/9VJcitfEUFkaz++T/h1o9sEsnh
Zz73M/Yr5KWXkUXJWAwzdIfnMJ/6Wh15r/P43h5BRm0A4qAq1Ur8KF2SOS7/TJgn
Da71iHIvUx7tkj/SQvNPlyXGj1kuyLgd3UjgBybgZwWkUPbShZPIjfj8uclybaZG
ZMHuF1w24UBBLxDUAorYPW9ZYOIxdBIOBVkgZrcQMkjP91gMwz/eO7bLyraVMOgm
8ogO5ZG6lXMLOUpUfAXhver0utqH8pM39trv2os/BQ5iCnNXypkP2YjibPgXlKv/
/+9bbA/FIorVwLAuZHQBCQsKkBmyVKsfY+hF/HWq6RLTxG9Sz/KQAu2+H5b8KLWf
8MGj8PONKzvUaaSJG2TWsBxYtTKYJ39z/5UjFdfJhab83rdGBKaoU2wVIUyXQBC5
Hscxr7bztQ2zDrVSP7TGpWptAeQyV4yd6SwKHeKVk5W+ggJSTh167gwgWcsYxXwD
F3ZSAjdcNSDfoRyHMo+xyUP+6zbTeUMoCAFZcnCrTvsNH3qOKmJCsCkJtL7dAB+1
x7/CUrXRhoaje3Q66p5ESVdtA+m1CgygqtyGwkyKTIO8VR450enX/r/QK+iFJtpK
z/ZGadH4a5akGxARlYWY/vN4wosVzN8ThPXMmOOZk+wjfBf/pqD5lgwu8NmcqvQR
9OmqIFRRXGx8yeVEBTY0iob20ULgSGZvIfFyg+7dUd5TrF4FGQvsJqdoyLNb/otD
k3vlcJGFVM8/HgWU29ADw05ScCOPKGUoRPrusbQN4r0bFLoAgSNXVOhK96oTE2ft
ppu2XrVIyvqJCb4xP6QRzGVl26LGMykVdX8lT1LdEBvRO9A5YryL4kfgn5vqlR+P
xQRTIgJCoxM1MsKf7VuMCCPzPJOdFlzh57jOWMc8R1pekJi5jyvBVS/kLd7h6Skn
xMpV27XBY0WY4HMVB5662E7xEryuGNr6twCuKjUUh75mg2R7sARdOAf3jsq5xzfi
rzA0mZrxYLUT+2IkWtyU02uWI6JkUjfOFY/QTCYcocLzxuB3fByoJ59Ma3Sm9cdw
c6ZxWLcYV2QFo1wt48SjhI4QxvkI1xooAVl9Ys5khTCnlktSi26iPZb/qA9dRz+s
/oRIiW8xjIJsEZGyMiaXYzUw+HINaNS+6xe5G+RQJlJonZGqFUGlwu6ToUxhjE3/
okMnLJGWxwavGZc+DbMris5FSh4QwMMPPPvE0+jc8anMBt1SrNNtfPT5oPqGAznJ
LgNDg3oF12aGv6tIc7Qywh9ltVrdC/MrgSUqGEZw641jLWjoURp4rlO0Lgpsz+pt
hyB3G3FozMcXHIs8pxdP7y2L88GIA5B+LxfsB3Cwb5GCM6sRhDgDgZRJGrOv8LyR
sNrd4WJZM/KmK18iBS7wngvtqfGa3s5OkzTr25nJpIbAncWgSjc95IxxNHHipJvi
t5hjFrxkFR2niRLTV4pAV5JVQtUoL5S6YknVPwoBd5e9fn4hRzH+DIyotZwBwZkT
LueixA7VPYRyyIPkAHRzJiz9hQX2jzHQEzvl+Oq8V9qHKpHHH6jhTBA+ekj9b1Fa
+cnnvxMB0Uy4OBGLJ6eQnZ2aMpLNU7H0JQ6K7sdn10OBIHtMI9i48/xb+zZwG1Wh
kogPpY8qoCENTOt6RLM4RXzqrvufdAGFM40Z/JMg9EUhUo1UKJMYPNiUEppfMC73
H4rXucwdBSpS59kdFxHFQBvA/8OJwxZ3TrilpaWZ/XHMJ4L0v4iT9t0uSfVBXVKl
6ldpTwfZSjvHs7VHqw+GbchpUEtMjyq9cu6ajlMobbLENnpPNvYM+bW97gq90mRy
4tmVm3MIFpdEy9MiiiBCTXs6iRUTrvx8a8NCq0TqBRoK19QSPgKQZdFwdI7pxTPN
/QPrGdsZKtf72jv9LOL26oIBNtkBveBSkg6KhgyDPcZS1/aiLTTdJFkSg8LtOWq/
acUwE1tSD3LKLEpqrN5FADalP67+yP/p0gSxK1vb6ZjBmDnTt7zS3EfqIsxn7/sj
sMmb4je5ugennJ4xu0qukO6ETbOV+9s9ld78v8RgaKjxEYoxJyNsot6SN48uRTnj
9XudbO1Q8roV6hGN/S/CY8qzZrioFsweoUlT2g4PjA1caP+dsZGjEdNZm+srLvDq
HhyURrBqx0fZQGXpW+N/1G+c/7ZTxgiBcVG8AiRnDXHbzbVu5HW/ntKCkOZ8oODq
2jEptrKYasXbBtrD1ifYtF3i86+/3C5dtAtD3d6Tu/sFy9Z5ZwYwpCok+fEx9bi3
GbdMB7w7+N5yJURkEckgVMd70DEGdGQ8Mvgydj5Cmn/jzrD5mIHO8jXkM8SQBUt9
pDQq8DpHWe1iimGxkpQthnpooZxKHtRh/gztzrEVRiORl2rtZPm0ANnrvUkvN2WJ
g46raGkO8bz1icBxm5TXSCQrVZuOwN6Zxq16So6wm+wTOh70DgTzGMQCfXYcBabd
v5NKZkzo0NJRRugSi9Ez3TdsN04wnyuC8XXDLj1uf8PQBD7vrEpvYAurT80inLid
5yKXpo7tb77o4ZQKLshXDSvvriq0SY8s2KfAMCi5uiraCFK5alCCkbGyzquiv8MY
H7ISuYeB5U8Kcs2vjxY2DaRszAwJL4V021JoFlkbj/5txbzZbDQdYm6sfk9joMzu
/yEm9Zju5lOrhjWH/ARFe98/RzuKhdGAmleERg3saSFd0bRtMMB/RqNDTSsYSX1p
Y3zFYTS2ORVtfH62Cxy4C5ZooP9mAFdyHh4Mz0ikChB9H/nK61Z9KtWoY4wv3jxh
NTwSMMmd/8p5xnw6+BGJUG8ZOaONE23d0aNnZG2/+YKngkDHoh8qR1zI9ZzDtLMq
eVXV4+NrHKncU2I6hzJXb6C6ezsnswOqKsdqDjnP/2gIepNZQRYfLt+bFN6pcJ5p
/FhbK3e6pkWlFYNvPWDw7185OCcvhlH2D8gCN0rj5L/JN6pTxd3zr+fW4BO4+yag
zEJJOU8Egw9dKbbRo4dDywD+A4Kc5z42HFwvUdoLqBkyN8Iqz9lgRfC33i6TpKln
4XCxw3p0z94kKVhMNTnST7ZB5wDklgkeEIJvINlMs83gNl9a+CKdsSMXoVbiHRY/
F9gAwrbzaDqpJJfCz0zwkUoUZL43Ee9iXytquL/uITJ03Nrb/qW2wV5EcKfKivyi
RydMCZjnbVcOaSq0aRJQpS/Efp1oiGlrvCN0mQo/PndtnIjNOieqLWTl2iK29qj5
rGCct0oOE3kYU+zf/j+IunBbvrsxenUReI0ptfoqCwhUmFdPTJNFTieCTa0NUYfS
zhE2CxJni9YmuLywnH23l28xjMJ9rr06F0nJ08fIMygYf7TmTPPYnnzE/U16EsR7
mCrrwaT/ojlj8jrDUuzHU/WznMF6SpSvRAfbrmrn66g6gmRS/1b+D9JfCSz+VYFi
d0omocvWT4r1uLCckveCusMXMyyM2rykvHq1qz7gJDYhJSVZZd81ZC+Mm04ZBENa
DDtYC3LNqtVTtJ/8UE+NKYSsqxIfMRf0DtjXNK9Gk1UDWlMQcwTHEjkMjQmiSZDd
AYRa/djaoSLo1llNJgLBXMOekZf3/l4fWRnZpWtRXjPNrdzS/wHYqJM/DzsbAc5A
NhTodzTD2DipfTo2bF2RJWIRZfDXs/EoDDRjLuxtobdFIcKoNhiNrDwnJGGh6P3G
aXHH29q3mKyvhHYX7K1T9O6tzfkCaiM2ZeT2DOGwvS7IydfQBevB9jh9XLcdX5wA
z/HY/iOPgg4WV6T8ZPQGnUsQEkLbOIOQMx0VeUZKt70BypfdLXgl7rlUW322TNlx
KUDHfMUfiR5W/+LpYaLais0tG9dDXgZZHPHsRc5RZi+3g7ZAlXz7/tKh7n9U/Ihq
BBeW9X+dkfM+OTMKcaJOeZorSjfiqBSWg/yEDh/AE2st/QVsJbmGVHmczJAF3ZqE
GRCcd49T29XDSBlfmjNUHaSuRe0Mi9k8+k7kobQTQ3VhnRfdsJ+ZDMAzH9KTCSVN
ptYhfbLrOzBlgt45J88HAil2czSsXAKT4tl3rpdH2q8bPpDiP22B95Uljpr9jQQj
I2Ca0wyb9DnvOqtZxTx7WjCCj0SPsXXHvGccxU3Q+rDqb/0IESCFBMVR9xiicIgX
Vj/puG6VBqf2ekDlUsRHXFcDb9NSGM9wLZESzdZg0o93cxgpBcb1rZaXwmKkArgW
W9ZJRzCqUQ7o44X6PiHI8E/tbWbtcXSGhQqM8sVu2iMU7Z+Plouqs3qdYDODGUdQ
kVt9T83w2UVNu1ZGOD70BumSZrpxsxQ7deSPFviTz7RsGKhtV0nvM+v8BoGS9zGu
PYQKG7wGU0NcFGvJkoArasZphINOM1/PQFUekK34vBhq8v3UH0y2qlEolCa2J3NA
A0fJoeM51QD5rfjIz/gi+b3lbjqsh8fGI4i/o7KcNoN4ZN6WkJuzKNvtXO7RSBsN
SsiRft4FAY0HSp9qPErMQWw5MBMeGoMoeLtwM2lfRRQw+bCX8o3DXzNe/c6YTW5K
UMaWcdsCAbDdbwoSgmwIJfj9SE2lYzGd6IU6IR4mDi0mgjjN+n33TJCXDGBKuI+Z
eWq82r52BV2y11onrwF2HZWvaUlmr5f3pI/zr5kXxzhV9NF/pdqpMkyyqIeeCkVl
WPvoyedDmySx8oBtHfZR3aldLNm7P9cC7LGXoywMiEobNFn14fpBzcVSM3rd+1SG
UbTHlFAk8LK1RXKo1Oqwa/iSrpSyBLJYkc9iZOxyLKTyOIzdoK5FElXQu0z+4Wk9
9AtWmuQ5QRd3lR1LKuTgysNxBdj7ld7EMhkyxEYlZUxIiJrQz8xMl3X3Yrwv61GT
enFyKkO9oDiclQTuPJTakndMvTxu8HKEn9iWnzpnYJlTNclspF2ENJEtc5RC02xH
nY9zLDjD8f5tHT7DsM+5hJO/4nlx6ZPyjVL15bJHvJOlVZU0qwftr4Aw9jxSWIvM
Td2fpGNnsK3dLbUoMg1R4EvMGFAwP5Wv+42/JpfHfbtr3HGj7KPqBTf0BsAQg3Qa
4u4v/syqknmfBSVOwbvJI8O8NmoOtT175y4odRIH64fVwNlfU//E6i0odDfoxFJT
2sko/XNpspqic/IenzIEBM7i2n3v7Mj0gsqR86bKHpr24LTj5OOZOV30I4waun2T
M+2UoDzROgkbhFRif5Js8Jo39Ei/walAhb31csERG9CTJT2tR0vic1+bk5XNaOrg
nmMAlG2xXTaI9OlrpJQggX+EFkFzaIMbM/aKYab075pf5iqWRXMjiLHA07JAsSrb
qCJAkVvvBsG9gN2EZuFPdXaS9RRdg/mQR7iTkD8wn/ifQCeO3G2Q4OMY6UXMgv0M
ZprdnmwYNQZj131h+vBkT6pNh0059km7U1qkrrnOimN7ZDTzL9Kn01DnSImu60mJ
mmxnyEJILLGW7qIHZGiREN7uw5wQqEj91I73jqVaJUWjCDsmRv1xji9UTnggQpJD
fmaPXw6pHCPBplR8hB+ZmLBXX0muYbTVqIB2cB2uN/WeKNFvs8r3iqbiJAZskQdd
G+vmCzsC6qSU2C2vVF/mo19AM4Gry9CBL46uKik9G+UVy29LF4MpPF+VVbSocW4N
w+tt/rjB1KwvSeR0Niyo1ygckSe3g/SlMECXvrkCLxDzsPFCS1TJhQONT5woMVUk
ydyGo8gKdp0aAJ3ZbrlPZ3e/63kvlLyqZUSa1BavvGjghP6sIGGjOxlC2HEtFzrf
3eYjWLzuu0Ua20R0g0qXF74mAAZqjjlUqBlkxASeHYL3CbhmGH1ehyzmxfhnXD+T
saTdp4uCG1hRcixXvczeVz95TgKiLmILI8Fs2HzftC1nO9A0xJhsRsExtW2o0N6G
xvl222+A6kqhfmFOi0abZQS9iGcsmeWkMAMj7WY1pxEnv31nI/Ub+qvgI8O0FH4z
i9507mh9vXmKvbeYcbpZMfDErlcH4d4S67xB/0yvAOtOOBcL3C1hhie3AXiEGBDa
QPJEJpvoJNXVTRQS8IJAbhUuRo+wr2zZCApuS2crabtAMQtw1LKNl857dQitmLvM
01uEUlmgO7IVR1QJ3OKLSqn35HGSA33tEbVNOJZHNfiQGMxE/isvniusgcBufHVA
WfPkAFZPZmVS+PkBKox7Qg7lsGAW2PPegZ9buAVIEAWx03QgkP1WAk3RUTqW81/i
8A5xTkVctBanUnaTBIx5Z2F1rAynf1lagKOXuA8ueOPovCroj0XN20ZFrpYidbBJ
fEu8WoFC7mgEhH7VBqrwexwm2qFo2Tct8MXp21JctGLkPESClECAJqsx5uHeiStt
gWx+U9eFIba0M1JYY4a9qQlRq4AGDb7cEJJgu+7syYmTr32PQJ+fmZzH0z8cOL7u
25NklZd6KJWh9MvgOx2pr+p7NKi7y7UX6qm6IOSM1Zh3DDR2kEYt3Afg51DfhM7e
EKDUFu13rS8P/iEWCMIeHdku/5QU2D0sBWomIxXNwD9xq3GivSWDGhdtZ8qCqG9B
4i9opD6IfoNdQZQcN4kN+qMwR7j1nQ3phbppRif/6xFOwuYkBlHfGGLIRIa4Gw94
6S0SFpj8MJxvIpXyr28pQOBT0HVvNIr1NhmgOmRcoLCeLfplMduVg3JpzJN+HNAv
2Tg0gLkPchFeOUEIIvKbreA/Gb8AVMSpZY7I9DQAkEgQg4zsAdZpxO0oE/9aT8D9
cl1HFFN/D55OHtXmsRmvKEvR5sE6YqEjgSdndZj12SiSUde0nliSZfjv3qghCFWC
8PoM2jloKRXWyoopdZ+cnh7jfn+HUvxz+3DpmsnCLk8Ui0c4JPCDpKU1et1ZcvUE
XhJH04rEXNv98HkzSJy2wdTps1yZnjvPkelqXe81vWhLvW+zzyPvbTGpYP4kUh2G
1o78fj0qGn7mICj1n05YDSMPtbqepjL2xO6icWzowFE5IwDMRIc1dKxuxrghBIxK
Ehr2zl3gEpSArkscXfpiE87X71a7MbhlPWjJLIjwPA9ro03hdD1UPVYvrui6asSb
VIjTRfg0jkAD12b+Ar6kGZWFK1N1zoK/KUX7b9iWyW7I5uRs/y4tCAKz7WfuEcEt
ZHTKsCZ6zEM3ra2pV5acGyLbiP/ptEbDKvIIbQWBVzRxXRpH9d3y1xJ6NM9OzcK9
Z9FiEvJGfTV+89O01gKqI86XKqYoB/2a8uT0oqNMMF+eT0TgZy6ahld5fKi7u11j
wZDZNiCCkKk/DgQ8lkXsP9qPl3id0NXXnJoRti3P1td0K8JghCp69uFrlDaHN30F
XbvIJDcmZzxDInOoXwqcbCz/BiB6hst2VJyOwSdHMBvbwYy5/J+G/uIDFb5rHYGa
sxQxzRXUK+ZYUFr5QiE0HlLK4Ol6BcBOL7t4/7ezdAtIhL1Xa9alX/L60/DCujwq
oHgNuF5ooZGvDq8wJc2tYku5mRPtNFs7h5GzIhd6jhgLUl2iabN72RVlUMW6VoKY
6DaurHoUGcwCQUlCeQ7Ho7eqzgTepcBMCysemrnG5BQqu/0MyPBqcfE1JwOSIWzT
WfaS6S4gWuGnWEDkz/raGSsosjbm8raFmUorbwTZE70NmEdpZ5FHePKJ/a8emxrv
0uXY+G5AtQqyfYyW+3eenbSHBmNnemGyzgoRsaqfD7jbHH/2ahPuTZNHZPY70Hzx
htLMqX3GfrAnyBsCWDzFvxg6aBVbHnJg1lFUNc0ZmfFt2d/A8BnxNr0avvlTfp55
Npf1EsVX2yCnRjD30zH36ia2oYA50yTh2hQSK0AR6CDeEjfc4SdfOOGhxXW5uZGE
Xqz+Dxv2+AYMb90+WoKHaI7NAEQ9KQrMS/8pKQstfOLxatwHcr3htJ+zmVO6i2sL
7OuSwkmk0m1XJp6kKG1W7vZANrjo0c5/nVrmcxd8LTKVd+UzWRM21t9UCAnLNmrT
93Ly1KpxpLtzpSneDMHHBOKt7xTUHzErcorecb2NKYvy3g80xjq57vCSo5fmjk9F
UhFI+hjITphcN/jyzieeieIHC7PgOgEByHXb+RPghN9vV87hNcj9DBoK8odq05ik
+PyzdrDr1YfPLxoi9mwfiFbd1e/5xyfPAOjlZt7wrONecKqO66D9IZ5mk6hT+bPB
4YTMAm3U2R00tSWvLPnneJC/GsJwjCU3pNdXYLe2VA2leDZvs2XcmaVlb7WQ6ZFl
kyGRQxOSnVNfCcaNEuUgqnIOXPvZFSkSkpfH0RZNB488gUN2L0gV5HobpqEZUCEK
UwqMmkXjQpiixweNyp+hCzxYREjPcJpGugndz6ZsNUjWvlAxX5SXgMCJLb2/5Wcx
6Ozoua8rpVZBHAYZxTfCklWPcvOOSMt3jwWzHdAMv8sI0fUAzR/7KDQ6HCFl658g
ewP5OifrSXhShzJyDSKDFx8/scsdM8w5jyvTUI7FSvmSF76zWmjGC34DkdQvg3Sd
DWOLR/vhb5o9Kj06CwJ1DkJQ8/31FMtzs+Q0yrdeUfZHWYA8+3YNLwjQRPd78HAv
9rj2BsTF0xj/X6XKxqYPzRsivyxm2r+jCdNz9y/akPksQe+D2YPoBwskZykvQlRV
nuIzhgDiEUQHl8j10msOFn6bBTV10LNdIL347lAF+fMrmIJnfYLj199jJE/wDi4U
Ka1XvK3vMIT4qBuTWGiG8xW8VZnmd+wx3wbSLt/hPChLB5vzIk3Nnkwq4k58CUGC
FnY3vAIPVfytIhwlrHtf+kz1dZSGU9oGdUSESjMf61wSzvVKzlVnYaWdRWDYt1dz
3ObFs8PcpjJw+95nlgzMaxKa1h0JdMaVH30Y6p9710nCmI5FEgDglUXLmp9fmTqd
Ob3v1WKd0zgdlpWqyG9AHa7jyY6N3SkIH5G3ioeBIHoDvnrsdMq0fYI200G45p7x
rklLtyUGjpKA+qF8ogCbeWUQQYWona8A5RhB5TxMKIGC+/FxWXsFkhgyF/IY8zkp
PHJmH8uD+G77rZtnNvsqCs+eP/UCSen47Kml6yfDWBZL1zgLA5JafyLiTOP8JiMf
Rr1aIRtV33lDQvlk5AY023ZnMvItGm9P6s4NNf9ztClgM+4G1WLjzmAFycSBESZa
JDOzAz/iVPPbMuC4kohZHLtKSjF3EkhCxxoc189ECMIedYIyMot8nf91DR8K+CQW
87QQK69RvvXmLz8/wzyvaWc7T2RK4GEQNo0BP2kz0Kr55+0/gjb25WIOyR39WD4b
RTqDb2sL+XErN0g2GH0i+lBUgD7iMhpA07oWgq1Vnu/jFRX8DigzU+gMrBIBK7Br
UgGW/PgV34sFW7i8zt6Vnq8UQLzKNxC5nsSllpR6k7KEkSe+6NBUQtSGalipaeux
ew1Sg28wDDnIv5Ql6B4AHyq9cEOzAoqXdNfzHKBAIcBknkS3/3E+dLzvjRZgkAG0
RBLFPm2ulOGScj6XjcYdSgxcgIPbW0TOCUpmJswxvRgNvepAa/gCub4s/L9gk36m
3QEJpqzZqZzZNftpIol3DGg6BuQ0pvx8nnZ2vY0YRot3MqVtmf1m7XDAQHyq5D8j
DclrKThGrurjuc7V1L2lZfo6vrifxGj48z0mHIU6/37HQY5x4YhSP9jenm5Xehud
CXXxs8/qS2Rs/DHvaKRDWWlgqc3aOcWzp9Cpu/CMEcqWMQF0T+xXk9ReJB44PJws
sT6lpQ3dO/DuYfAuQbgn2+Kmo61QnJ4/LNRBzuvPTJV71lQ+G8F/p4lYoDTORwb7
Rbm/Xh/BRFj/we+NYFb/Krp9mVYvuj7dvkjWyAemjoIi+7lBc3Gy6UeTgXV+xsET
0CFivy0Xhd4ndzTvp9lSEIUb685AE0DLbLUuZE0VqJWYNfsfycb+Nkxk3Q80yemY
9/PcSQgcNl22KlQ3eIcaIljGlg3GXVIZ1r/JSkOv6yQ2tzrEkGeDiiYAn+07Om6u
bOXrnfO7ASXe3173mYUkE23NW2pXEshXSNYnKp8N8c9P6/8U0F8fUVD53F/ezQKU
HY7I6+N1L+vD1E4r65l4QBuYMBGuNU3G3urOOPCOgoz5woROMThvuO0rsHxibgn8
WTIKEgVn1r902Htptp6j7c7qVX+UzdTz/X8ow6HJUYLJ9TGQGpFCfe2u/g11qdps
NO4JHrADYfHwxux6kIuJJwv4wWdTBZkJLiKQ0Ab9Q1/aEvO2jtcDZ5+MNuehTSbx
t12scHuQZDosWI6j0dFY7b2Vd+c7PBN0esHQLu2lvSx317sCf81MqKhfwr1r+qDR
n1k7IN48XsRLY8bqCAWZJ3pT6p6g4P8wvQ3419DY2MWGBJQXU61LHW0+rr0obutx
9hlWQ6zIMUGhZ7Exagh93F4kUaLRVKK75J7ypT4OKy8nmJSHXPfGdDeJXp594X1B
mEs01n66V4164R+HKXupYdIGfoUEvTr3F7TDtJUMOObgd9BMBwAYOlwd56lIU6d8
SPIdJFgQiLHrNGHe/qf/ZEx5CQHVzR1EeTe1wa4yDq1AVuj/0Ghczccm1MbSz4yy
tlxYuEZorsUHKoKonVQs9NjBvKkpK/KF38JlTHz6FxKb/4gRVLyyHckpZRaBHVBI
AlWqKG7XA5wec+b0I5QoTYlNLxFOpYOieJkp8IStxyHis0UxsTdB9JkXFWtA2P5i
JiYnYLWkd9G8HgQ6SZu8amoBZGeKftT4p8sN5QIrG07FGKsOqO9jAgEIpIAknKGr
rWQ0+WxL8KemqJIiAxBrahgoNAYwnw1SN2cRoOYZiOLaR2oJ3LMiYC5PJ1UjoKcS
pX0ZO6ji7xGa+bxj3h3osCvh6VQRJigibCAvJuYd7rmWUAUPRX7pCy2ZwC1WC0H3
GguqYRvxbPZnJ4k9XCemCt01DE9liA55C5+VLyCZ01DYs3GOQjmlzAwJE7vc6LGe
RueAjDZu7JfcJSivN8ShtRIc99TG5+9/pcu0UTctWNH0UnyTxaH1swijOOxnYHll
PNvH4AIYCeWk5jGVS8p9b7qrRqVkmezRq8i+BNaOmFeGwfOElMKPgNyjnOD6GWLT
94BA4SJjRNIJStHDaMq4uDMD/cHtMe1N6qUF43t2DgHoPtYFYc/Tz1SWloByb7vY
eBflH9yCErWyMhNfLz6Z65wJlWaw20QTphF86y7cNli8wzENXWTZKLTS4X9X34Ce
razVhzZnNgKAzlPnu+7YPvZH/Ompm+zB3lTmSNyWd1eQ1RZ2mJ7kLmvKDkfU51A5
xhbMMj2mNkJUe3iFppo2+d1Sh+HAjjxsbV5CZs+Z+d80xAgvb+5wE0N8GSydfa2c
ZMX7XZ4tKW8umZSQ5Xd1n6frQtvvS5IpmPY2cjakNHsqvVN0HCNlgw4VgoQ91pQx
aTRzFXJgNOLsnJTGIFrpRiwsN+lkaw5CBYOnjbw9l32MDykS2gj10k0PTysIYdha
cwosoYP5u8iE+5IK4eHZt3SyxSRJZ+dsOX33a52OLtDCswnP1tAOJOlBDdryJTJt
CKPL1Gt6+I00wzgAkhfsqMfsjOqIAL35fol1+lemnpTBTZMeU11uM6s80V0x/PoJ
6WCkHyedmUKpUx3RN543rp8fDWofvOH6wdDcNiLcBr3n3LKjkjt1tvycQF41QL84
Id1RBPCiHYsg4CXvQ4ipRfVrGi9zcE8hw00WGez7tChNG1c3tIS0phTKOtCKjqo5
BsmF+pCgPH5fgSVIGtN4BW9Z2FjIa0WeQ8L+BV3imjsLtmzWKi2kCMib7AdE0WGN
QO65X7EiARF8F29uxGC6ZKgdujUtDZu2vHOgYgYVvdBUnnT7gWZjBJrrt+jCrgBN
lsYcCIw1aQsx+3kWeq07FmUebb19Trl6NUdY8ny+hhgzWChQ85C1bM4mhkHmwxz/
AVj0/EAx4GJSv6q7fFJmTF/KQPGTKzvcftsksY0PUQjiblPRllI2ErCqny/OWj+p
E/f3SzV9guoefdGpo7/xrHt4BdzvaP/5Iq366LPETyrd9EU2YpKQVFKMrwn17cG/
bY79V8nx/1r8e5ZNVIzr2FwHGMU2uVNqInC8vOTCokfdZpJ5dTHg7K5g+/Yef43d
jK7MhoSZscrPt9WUhBpSYYrE9+fPRodDOKW976V3oE48VbJE53A92fS6Q8XjnxDt
GBj2A6BgPEO8XFgex35d3BoJHcSuz0L1KbP8beOjDDKJZ5VGFY32kqADbALNh+1Z
CfewZ2x0pVsfBCb+P9W5ALWlXdVcnwDxF6oTzbBmV4Vj09x/YSK8FpbU469BDnDD
r97ze9rqR53HhJ4+/95o9O0CcXTcjgFElBuPYUdrgTSww44WfPvlpx9Koux6SHyw
XzRh2avIYaKJqHufC1IQsrlG30/vQFshrYmgK0iinN/Fy3g/e9wxdafSHeSiyVR4
wW1jR/3VjcaXlICsWPrPMUWXZcoATohf/0k6XKsYVPmTFoVpJE5KueoRQaGdUXQ/
BNseateyuZ8DnkiU6MvLWoV3OJ5a8xGsipMg7vBRcruqp0g3oyhuWcOxn28EBPSg
eGnqSmm0YH6YQiNF1GTawbAuqiP7a99iImj7/OKsoFgG49KMAEM5g+c5nKy4A7O1
4B+IXu36wjqB1mKjhk1uVKCmFlLYqJ2o/1+ySpwo0PzJrR10V1V5/dEVMk+W1dPJ
bqloAxLbBiXPkeX4V3T8jD09uKXcPAGf8QVxocASV8pWQl5YyNrrkngRGa+S5MsI
/bBthNn3ihotfuFG2lR4bSBtN7DS9boVoA9IjhD4bO+jwWUsgISNolZWsdE52UI0
NCjOutG/pcYUorgIph1DjrMfpixBZpzbwTUOOeD82DE5D8yLuzMjF0Pd3zpKLA6R
EnwTv8/ZaK3SR17BPZOYPeNkxWs7BhMuIEsIOPu9bXSy0/Lcflzb+cqycGl+4wAH
uRr+9nv9tObmJiBOOSnlYfsNAHxZY2fTbkB7066QPsxlC/7AhhgleB515S5aaDTr
JgReb8cuJPNwV+gW2Wc7ljDWszhh4VfaY2DQ24hVioT925ss1TFTws4K6RQkZMmR
BYGGeFtSLWw5/LyM0U4XvbNYpbcaZela2/Swy8KhUS5eiTWqU01/xAxIKAcPS3WN
JHQqTzmV2+FOVtWNl4bzQczDHQS3uf22+1i3RDn0lDU9dTL2Svqu5h4DsLHkqdo9
XVlKr6UTu3RQ8FzEAMDF+a4ZDWu8KbrZSMAiDlZhoyY55KE7zVrfpiYSmL3z7EP1
4XpAsi8m+1M+TrZn7mYifEfy05AqasugyiuCcXqMInNKVs7fJ470nYH4n8MntzpR
BfD/NMgeOWtWZqjd9hOvjab7m/A9GHIZBM1cAB+P0rCLzGIDut1QHAqtSAn6FVoS
uWAMZslj+bER49flcqaf7v539mqGMrZI8YxbEhxHTrMK7hEoa/d0xlla95ssBKAW
wsrYmQm+1aWjQcOhzdRQCGp79N+gTqwbDT2bmPe6Ue8FQVfkAA3rgPlKMmbDwmI1
s9Os3EuWhlDbFBDRHSel8YVhRP6nsVblgMNRrpTFEOunDMRkZyQDD2Od3kj01tQx
5b9sgZsje7mCH81vj1hsrtRkeQRXJAm2IDyd0390XXRhTmx0BCTpkqfUrRVTWdHc
xqloF0VR21bSmnoh+jtjxJ/7iMfsU/qT8lzfW2SaMmBDha+23g3+UWoSq7olIYkJ
I8bWizOOeGAq0LQsirjQ32LLraNQjEs3l45feTa5PYB6C1IliCD1pPQ6oYbHATr4
KzHuEPoXQHP5/shbh5K2GchijseK4/YkzaW8jXlmSni7B6PcwK+iPpVEsXAIZL7F
3illgWl0CeiD2sqm7yAEYFaPQW+Toh3i/AkXXd41l8dD6glCpZiC/YSnrpSzsyZp
FyedV5NFY4HmcwTRgRBtTBXn7knj9OHsETodIS07d02TeLVnQQ9SNxFyV3vomVxT
xDCOF6Rjw+B3TAnE16Q/6AdPaAx7KbucL998qVSf/nV6Lbz21YUQC0H0xquycVdw
h6nW5+HeTgdxQOb9M+mD4lsQPksVn6GzUX9+pm3X7tZsJUTcqntogRDRfSXxQwov
pgNRv1lTpA+Ogx02oH0mEQ7L8SSN/Z9dOZUnx4JK6npNuLYNZZbz/O6W8wN4gOFO
poDk5ly5bB8KOu+kvL9LQ+fzpisq2OBglgsnuG8uKP8EHkdRpcwGWSfLP8GKMxYm
N/fya5RvnqBcjFqNuNcSt+c2rSW93NhAQOFjgqK7oXJy2qHmBFPFV1YLtCaEn6IJ
cWzrtCCgNvysdyiCpwqlTl/QXiZoLdsHAZdE3QDxbV3WYFLBHYi2k4UdSpD0GnSx
jkvMzyNRLoewckZmTZHa4akXOdvXIYSEOVNtfR4UIlYDsOzmPn1TdvCSgAQbzfoP
gVqjTUspH0n6K90TTI4AAOdOBdy1Irzywb+jFgPeUcXe+St6mu0ZTl+TZHEbLn4K
Qzs0lQow1n7kOMdiKk0pJc8IFe2m+iUN3p1u2/cANGKdZmdRs5S7nnsMr+yAN8Ey
r/lLNavXVPrcTzmvj1oKn8OmVFhqIgvTFFsew+VD+lmtXkZLqJy9a4tYNQx/v2EV
Q6K+g4nUEYG7RErYBZG6/ZhFXJ1YngAtOtep38zvHbbBQ7ys087uPVplRrEESOz6
V8vsD3yap4B6QEA+z9SwmLb21ponfF2IWmUnCpmYZh8JYgceY9BrtNUWayd8toHz
+/3ERB9YkdevBkJTlCnokkVvHKAS3NC7iK5fQkS1BRVw+aH6o4107GST5HdCvz4G
a/56YO2bFSjrjK/nS4BpkKvpMvI2zMzNZAejiNkpgv7e4imj61mXhvyxlMfR05aE
IHaE3P7Q1/plNjrBCQily1UaMPGtBYQdGR0dOL5ha/svB8F7hRVtRVqNCn/bvAWv
M1Hij02UxAu5Dx3eLGN6hr0SdBkfkNFrXXCHCqPcunSj3SwGli3GiM5p+fqVSXAJ
jee5G3aKBS7uW6eWK+eZAjJP2UzSCHZk5BQZ4k0sXpT9uRX9kVFnID+d1Kis9RtS
MbmXecirT4OSi97zHyn3sZ6VTq4di1ihM2cUdBJRjva9mvdYZutZndG2gGuFf4yU
08Br2eNzXMkotOYQqlKRISsQnY7s9V9XOZGRlOQ1L7QKXW9mVJptigxtDXEciPwz
hfe8c/gkrBAv+StDryX+W8ZkHrIuOVVmAWyT4UyUOL48GUoZNQCxpYee9qod1cTG
YWC+3DdaMrP0Q1TfAxhz+VnesXAYCVChDDW7FVjJ77CK8W96jU7xKDIrHNcz8MlX
VcwY0lFxxqx4f2JzixYM2bUIC5tY7wKBInKcR4KjYZuCqLFYodRxSTJnrZI/ePxT
NEjw53jbkqpU2965NYyXM8urn+YHZlspuaYN7m4z7CXx1L6tqcGB0r78xYkpmmcg
K3R9vnEQL83uh4zlbO4P2l9InHgwh354OCseDqrL/fINAvQIFVGIV99iQHvnjTgD
AarT0jOijRyMhJgJuOdXUAYFWaWvnH7Ko8fnDNyKn+mO9c0XuXk6MH2C3Sa7/y+Z
XAcUzdfgn5tpjHEeLUwpCBIDRzEOVFCA5877QAbUr/NeMbngiuLc5x+mASeNHWD3
LF541AFpXiIhTBdPq1H8zpxa+l3Rkws9fCCiMI6/UEh5t4i8wZrcI+exk2sROw8D
ftLdilRcjDCiwQcw7xRDAEH/lxXbGpSoRcz1XCzICcCRLYPS5jndpDU1cVzzmyAR
YBC9gXYXPjWDpmy+bUF5db6pvLW3aeOMnbzQ033cAuxJkYI/NpQu8XDr1eMbilBt
QLWgB71kIFA5ehWizUlX+pfExZeFY26HCHOpUCv2IgRlu0MKbQDCgGEn6WUj7PaX
iyqI7b+VVdE5mNK1yYPp+70Nc92kg0QYHp6WLUAHv6/hazGD85TMGnCN83ljCdHC
EdySuzD2F52ZX7UdpyaE/lAVtuAVjabQICQDUcw5jifllWjHqw2e7BXMhL9IuEq7
a2j8IfQRegmzLBa3m5ePDwIF8oI/Ly8tktrVLvv0H6tuH41NqsBR3IBFe0hqw5J1
IV91fxMR19LAZ+X1/1eZ7QUlImTYlb5swL4jp6KlhSVbCYaFxKAa62I819BKdEBR
db+i6qpZ58x56j8iiLccbAX0Ba6OPU/DIQudmHPGcqkm9lSwSGhGhTBBEP0k6qrB
7xEBw3q6ahvEmGSknLM6pe/pmSiUZJS+8dcPiSfQaaGEuN3hiSirE6Aj0RbhMAP1
Z93bp/swPSjDQ5gk92vBICnkfIjbqUKQaSgm0qMGaAlrUTC15X/IgLY1XumPEtol
EGbtcwpDS42R7OkUUPhN7XBVsnRCN/+SnzoAKBZdCwuMnP0wyD/fvYqn5JAeYTPj
JkdFPJux5BOv7jPTSUSY144zSB6e/c0G6joftnyv3i3VtqVJLmfFOrH6XlSfpGo/
BIJ6iYcMBjuUVhqbeWMR9RLCm1N9tTdnBLaV/ksFkEWtqvyldd6VHOkvym10a6EQ
uuYOtO1ApJD+Ew2dSG6XxkS2ZmOa1jbQRAlNAiRWbx045VoQEgQ44mAuPsbPDb3G
pgFj1XCXaYsIQwO6+Up6cnYgxbDSEdwKzBReX4OXAB8paKkyEYzdkLOPGNf+MxED
4F2ZbTFvoU1Fobxdukji66MzHHztmdSIW4eedfs37HX0QiBkogM8igD7lInopyfC
SVuuERrufbFqHF3Tob/mdc6en3atCXz7NlyiTa17Js5RA9gQ3POkjk0n9S2AutPu
n2d9+20BeciANti3dDmipqIQcDQuIYECvSTl74p5K+Dh+ERAwMhUWRosixNXZ9Tw
gFPz6wiDFQKjB8GGnd4yqZVqN0XdrQf/WL2zHhVJ81HIecfxrrglYVL6F7De5VmL
U0jrWyn3w5EIfxlkek7oyCTNhtsJJt2mw44rlUZC6kRxmuVDDOc8SbW2eXA3+fsc
E52xMmkjXUN7cTEYyPBmaQrh5WWwqLstVTwvwLWcjY5/r7Iz6R29EtZEeOwtsCck
cwBEmXp2mDDpXrMv3UF7wZs4cvVMDA/gHNz5haLUCtQ+872ncoI5dr++CZx7CNTe
wu+ayV/JWO9/T8OVbVuP0GMI3xMswodp9BOuSThz0jBN2QuY7uTSffkcCHTx3TTe
umgSgBLcDtUwrf/It4DzXzPVumvoRHM7fl+N6UVI32uSu8TnxK5kruDUtz+AhcjL
7BhESlhgTT8NHfC6+Op4tvZML2sj8Fqra+jOsrb/uMwz4fvSI2IZolKOChhtmwNw
NmUnRQ6mvAkWIP/qMcLRvcyXhmhP0BDim/Vh31Tc32nIu/rlk+eVkkRoJFVsFirN
688wFmbIEH0D62mUbdZB4MKfpnfBhHxoLsIkpt46ZNc8yRo/OW+NDOWwC2wfD4wZ
L6w8hyBY7/erYeOqwXLJjnsqpd6Yt0tDmDefaL83g4oOGo08UMDVIlWtnFPNh+69
fyIU/p0UpOLz6QAIeGXORku6vW51St7CY9cOyUCUXQRBcidDG5riKztvtuknvtrK
u7t7nj2nYG+yXtDfqbPvuWVh3Ik9LSlUSV1496siuXZPzXViAIjBG1oWl4xrHLcU
fzu/afTQ0fDvKs6uInYWXLFUnRo0hKjXP9RvJTt1TzUhBXmOeH6W6pQcgcEVfI0N
jSQ+aW3Fgd/IleeRSdEGrDMfglkKB26dB3aE40qJNrlEggcfxVHcc1kYn17/OG+F
YOP4H7+sZM+4crDedz0exE+/pDqzuz5GQG++0fPvvRQO1nW0E+8HOcXTElC++AAT
zwrx3LB0+fMIgfrsOdUuu8uPKJBTnqSBisYrDu+loGsT/owvlX5/FlkSVQjGWR0d
Cf6A9FZKjfxSLf4B4x8JzFE6nN+uZ6X71VUV44gL8suqLGNW+2n3JyWpYJgPCMF2
8S7hySO76R1Er0XkCHk4OQnBu0unfTnyE3F0t+hgz/RJoYprtPdCKA77YKaRuVuV
oqB9wwaquD3yJJvXX7Les/kmpgiYeXOPyvNSXUXjtcberldkfVF3jIMlghdNUCa/
QD7bnCAJkMuRorFoq1U2r/X98d2/VWSWLLMb14hINexn2TjiZb9zITWO+rVMRr6s
FwMQ7MaO2yfqZlCCGrEbiFryAd4TmXxHBs7PJIKVdkIWKf9Xb+0CwF/8/WwOXYlA
53OBzmF8gUkoKBTki7ly5IJVvPFbwqwaGncccKeT53QSjerDRXAxOMIWqzi/UNWQ
lIaITnS1ZuzCITmfIZs6ea/MA3HOxGl8frsE8ow4OnQKRZ68SaKURK5/RMjGkwKW
NoyujhcprU+P8YP0ZTia7t6qvI/u/1lVz94BKs3WeTsDhOV6kM/a9nAVQtj9rqZQ
iM+F6jlWO4wkbq8kS+x1MB8yLbmFltf5oh/CPrmV44kUeibrLrtjxUk9M5K97jBf
vYX2TJ1qussItzIwQmjwU7DAxtTu5EvQ6WORtA34RBZzhTsSn9/pJi0XFBn1d506
NpSgy7wGlhWbsvJc4PNZdnxMcKwGD4D6aVEAoa2n6GPlBiYoGyc6mYYoHk1r2RXm
G+dTi6FbZUaRDqwNXcr2skb/qoKhqHCgCvNZzssmZmHHiT028CzAdF8eJUERD38l
xzK+OCW/REsZ5eq8tzAz5jLEsrbR3ZJtdPlOFTy2JMvfS8PQXb/glyPim7OEnmcB
Lk+FgWcAvs9Xj4i381LGn9WgDnykrJmpuZ4sDq6K0Ma89xe+tG4/ZOg9ACb/1WSn
XnwE8V71WRIx3/Ot4JzyCgbMWVSvnlDUIIKgRNioLKboOD/25HgwXuyLQfssFay+
QqslI6S7ZraRrf/K1TWD7Tv8VWgbv1WaODIWtHjyZ5Bs9egdnlDAn3mC6uVlcIic
pzOJgXds8iTPtPfcHquiactFg4EcUwrdwUy/CBcM9yOsUZv9nEcCugbzQ3Y28i1f
6uDlJy2cZikjQMl5xA3H20xTrDywmJzrZdEqjBEyKllnhpTDx9IHhOcAXspj2n5e
GiDWGMRy0YuqI+fuRSjCLvhjvGAKenzdMrYykvrfLw4+3SoRwen24VxM1O5uvsKW
l+OGWQx/sP8+qqXSszzvAp2Nc0eHiRyO+j73EtgRCMHuj58Imo7TI5er+xxzUsPa
lD9WoaFMllbQ4nmLtAI5MUkKgHS7LihNLb1xc6WHSUGFpfpFqQ2vB0p9ZB1dysQU
hwfI6hpQH3WOtlR++qkAWbYXgTGu6rzt+/3iiRx8GaTAbk5+MmU5waH8I0VMvyjG
MaWw5nLeuKMY9dyb6kv7UAUo49G8p9nhEwJUWSw27C7uShFHNWy5SfbN7PUs6hCA
DLFQUQoRN4YWnLMW7ZEcIj14eVVPOH7GEinJnWwoavlHTXukJdDKle7jMkmp9CTI
va90+aIA6uUc9W1HNT94vspmfVsgF0A6HNbLCauVtQ1cW9PKtxx/Wp6bwS8IZyr+
+EXcplkjmFHD79Y8E+lAPAzVJ+axiTsaGNNI7v8oRbpp5/mC0pYlEYvXd6HvCwsR
vMveo5hQ8+XN8gYBfJy5uC2gTf4D9lC1KB9N9OddDcwuA3KRCwFWHILS+RJlF2lc
3JL1Tqo/qlnmesR56zHvpHMzpbaZ9Zwg9moe4vCzCsPxms5AAtmmTvt5LH6M/IQ2
GGmyuv42EBSf6n/Ng15IXc5vzOXpBJDDaOQAosk/KZEw2hgsfqziR+ueFBcQjUNn
SU3uhLXeRlaMqtGDzeV+wyb8UcGLj3nMElxDpi7wwa7LmCCWdLXc8sVH1sBaHhy+
pQnzIKgdDeVH6lfJqoeRKL/iU+qtxDx9FVNxq3Se9tGpP5Tm5tu4udvH4QEgVvt2
m99XZz7E3s9tLUOF6A7cVDsPxs8tXGr3Yq5bfIcHaTZg9lSdROP2bu+ftQV5znY3
I9aEcaokyWhyGGHSn8tgV0ihzNS9G4RdQP7TkFyWOpqqJKfhEYKjtEThumljP7zs
kqyozNWZtfcOXeJy5QGkZJpxbMIEcztfRR8rhGV3u8JLJNtXZNiQq/+wSBdcuE0H
TAAs3C8jRoy9bhf3MBEQxpaGKHpkgPMs+87lRv9WKRGmsln8T6xrtSOgfVxFQ6hr
EEgunyRQJzlLs7TDon/jDq8sitiM3y/y50xSaIs7HuNK5X/UkUm2FLhWEvsdXz10
+rWeqU2b/8cRtg6zjLK5NrbHlrITx/NYs/oGCu6+TzxCGEBLPox1dmHlixpoHfn+
dhtfIayy4Zh7ZuhW7JDmw6lWGV6TWjggTZTnD51f/4aiNNZ7dUklJ4uZvpN6NNEg
RDDpyFOjaPl0RXSaAhU8Z1rifFNZeJh2zpoUYyQntZaPdzA3yk5BTx8G6InUtfQK
j4yN5D1LN1qUfN+FXrWfrTVbP/aXS4NXKM8ouGK8ToRytVaMh8wvfAjtnbmfzWui
gWQKBckuUS1ykwN2HWM0qk3VwbOmlu7dnd+wyuTC+ryKB4/RoclrP0TLLcfRAWd8
cuLkVkP0jdOX5jiVdt8cRkI9YshsV1GgHxbOGi+mJ+cZyEx5tLsasBFfKWVkKEyC
8I8/SiFLgeXkIE5Ad22VULcmuJc0vx6Re5cNunyG/3wsUevhOofBZjrsd6VXpQof
x9MRHJ8X9ptTB7SXcNtMjJcbtrpEGW5Zp6GmEaDtHM2UVlQ6N3bifAabooG/WbUb
yZ3IfaGSZbRcHm7TKmef1PoI6eAkwWgBu/t6XFvWLTOaFM9hy4FErJ8myUOwsEdB
vijZQbhxpzjA3mEh61PC5gs3rMx7nb+0zBwnufcSeZ8UuN0rjkW916bl5nsL9q2h
htmxcpzXbcxP4affpG0ODW86p1D4N0tm1LtBCHUjbrvJBt2NUW2ujD09JEMRRskr
gapgjW7Bm3fjQsZp0y49zxgVwxWSq6E4FkCewQP9Li/iM6o2fPkErZMhmQP7HRW0
0hulNJhrJceLp+tIrRXh1GvzwlNWvreUa5OzlTQKHWDjGwjWpR5HRem+3h6Xm1rf
cTYNQjoP8hn+W3WOHWR3K/UO2QTxDyPfGX9G1w/wteDLFuxgU9R7dmSNG7EmbWlX
i0UCJsbkp6KclRhEo4PojJUDmuE7rLld6saNUznzSzUrMHQU9EctJJ+SKvRUDxSt
CKCOTW3hMSkOisBdbf8N87cJNFzB82GMV/ypVxBYN2zkSYrpDCDGw8xrpBns8Xnw
YYlgXkDlrky212YGR408Jp2ukJ5purKTNC1WtYe1xnNjqqbGYzNGgCfMqR5kGSkJ
ig7uJPbdeQekBP2uTCcVcrBpJPgIySiPUa6C+7vPZuX2hu/yIJdhw+PHTs1oFcBx
gjn2o5lcSnOWJdxfWyKf4PXsP3nd0KTAtKhLmpS4p80PlEAbaW7e7sRG01UMlbr3
Ee5W9qdFgawwf87NVeJDwHCVaxv7I3N1y+ZzDtZ8AHDPwUlXxU+9xR6DmI5EhY+3
Z9g4EMqRr7/BPJAEjV2CHep6O8ZS3/EZ/YpM2GWUIGOzbCyzODuQkwbb8Z8SMS6a
irw4DJ2e1AcYbcF1bmYk1mlksOzd7/kMsTliseuTxMHXI1RnX/PlKi4vl4I7dOa3
p6GBnO60qJrBBPfwHV9vK/n3eoMaSOlSXCjfzqS1VWtJ1RPA11wRvgTirI8ITP1B
YXoKZw7IoAd/Eoy28l7La6oabVBmXWGP2WWOlsmTbjF0iLIfuZ3884oEtsD7LtxT
F3bd4YQsFnXwHEmlxeBSjEKRGg/pdBSdYnp+2pMLTwbA5HrIG5hZiHZvGA2HeZ0q
9YivdkOnMoTapiwnrGs4Cl+PAkz+8l70PmvPv3cl1/3YAkAl0xd59zgk3ztP3If7
t7YlUmK2navkAXI3SwVMjPQp2sPwcWC3PbmG0+x63zPVEJytEKijsJwWZfq4aE/R
gXmM8Y2WJmRH4IRu7d2DWNXBsha2PUoMJk105mFEByGbVmfGXlXX2zRBNhh/33sk
pRKsXmXogHSTtABbSirbQXCygAi6hhzNKDmX7L9GpxeYgFpsHqWZb3D3wqIXFiiB
wL13q6Fk+8HKrkNkk2DQrVnQqi3F0A/XaaS5ytkCB28ReO9QmOpK7P/cvyHM/K88
8mpcHuzqpNX6DNQNwaHTYA8pkNvrNX3e7fmio40Z/8+iTB2mMlHCGjdRyKkOmjJ7
AVeNiBwdJ08AThCPnL+c5P2dZHsO4JBe3Mi3yBEqPTIAXdkXWEyWYR++hFRUDc9W
9tCiIC+0VvxUmI6CMFVZCHrokNL8i3kSrKWXJLyaaHHWH9FLST4JHwW5YpcxyhwD
8HSqVgzMWx0G4quA7odkMBuCPVRAvZepyKw5CxA5y5SfqzKjsoEWYShBmllQ0tPn
Y91Txe5lIFnR0YfZyuHX3y/NXrvNTF75Gq3qV22NX3/yVipW2Zg6Vkyvfxr/lQsg
If4IjztOY+YOLaTOVn0mPmAfr70YedPLb9/AAegi7LkKdvx2zZRGENOY55gDNioY
AqIyXNEBXotE+1L74653CI4ebLHoX91g2uBzOzcArAgaiwn5cbuE1ZsaW5yM8e7M
sQ9H7Um1jaPNJQOHh6ascPxaSCLEaX/40OBo672UQl9z7U/c5RF6QKu6rJVRDHov
sIq5utjJsE0wOKQrGe/2QJEDoF64yz35b8JYz/2IGnqpgYhHlYpVIweQKs25RLX8
u3eQrgv2qSKHtuJ3OJJ+7EDQsUxbBqyFtntSGOP3lWJ+IH6Mwn5QIJvo/mUUXqgE
mamVaYBI422jz6+uAMnScvYcsbk9xdPbvVtZDYALX/Rz5DSullLYXXSJLaeXoa9Y
igexe4FkprxPyBRmFs27w9UMSMyymWG+iimcEY6k8uEU0PO6DWl4NEGuCQk7rtZd
gA5FFFpiajzndACEZ5642f6573MZBVMyOB9ZbTZQpZIPx/nDMY55cJ1DMp8j7tEf
70to0EXcIe7nFKEEQFhwyd11Pfw6jNBT1nnUvIWfSwYYCPYaw86HO81M+KpEVzVs
7XotZjFsmOH4Vb0WX1Rn9QClcxeHyiuB+G8pdo/XcJVsB0Mw+Alnc0YiZ0NRAxrs
qDdLBmGgwiC+/lo+sAhWo4ElBnp0BCfLHNOFTZ8DJmeeCxQlPEHK9zL1u73RieaU
4vVwNwFimP+X9sK5tMi7cZCriMTPKKk/ha9hnkB4ARV9NlwxuQSc7JnwgBjlKheM
9yxaKurg8a4ER+1uhmHf1gQvOm4kTvIWMqoTwyYcy7qHP37sMV7hLrfZUxUa8SeP
8rXTMVYS7h4c5nQ9dYlTUzY5l9oHPjK0oKkqStfMwyvt5z/X4TMlllE2Vf0Pt5SM
lyr29Ekvscrc+DY0DzuIFvgznN5czl1uyBaXPiFdsD5VMyInxfVpXURJdgtrBtIK
+pCNAfxZxY+qxd8fbQEB4Kw3WBEhD+F8b3ka0oqAPqXW18Si/GTbGak/yI5m4Npv
Vii0EeoWIbiyzCI5KVXdBzlzlIwuaHvOg7s7owbViP4z/kx1V1Tr8br0Ylp2H0aP
3+2GycomvWA9xtSbmYk9xGkSu4omSDlvVHjfdBP9jCy04RRaguwIVszAk0HLSWHX
4K+U25hP8OplkkFFDoPLcFU4lqrM1gAe8XmAq6/n1EqP59mWRwsuFRt+XPHTNOex
b56Ap4+ssaV+dLCjxA515P0XpOMWhHtScm2uNEelPtQgXLnd2+VIKvpVwBEhxmXA
ShtNCQoH5oJye2qRe8G+9M8SRCY7HGTySnOHvzF0Ti6hWCsr/J8uDSDCtFpGgtW/
J5SnX8sJXJlHbatjralhv+LR8i3ls6rE1K6dNYn7idy9OtocZhcXSM0/hIYm6Zkh
hSiBWpJr5UW6u+BljOcnwc0i63maCAXAGU3CObD5QY9co0ydfh/4B8vDrApvXhZs
FkA/zLLrhJs7Wt4l1FqbOFYrOHfM7G0f2SXddmNlSXpeS+1zVmfwWxIb5EMEnjD8
OfL3hPhowj0TtR6ZPb2h6D/0pVnYAZW2uBcQcdcXo4zbnTJPyPzo8JUx9voYrWYv
OPMzqLykgdfCftGT0lHZ/n+jqSRcVKSC1KihHAVTexGceBZztSp+k2EDJ4Kuc7ID
o7p3N5+mnjPAszSVFPMsDT1O9o5joRx98sSb3K8ZYwlGCXzkWlpJENp2bRA7vSZA
yiClpMYYWwlzp9IFVZ6MDzLAG4/pyJyE6d9rPOHVMC/1MoQAi2BDNrhKuUrnD8KB
dfYdyUAAzmkt2UqZMf1EkIcS/9msUVvmu7QTFrlibssEuW/Q+jJKGWsbBDQ4nZA4
bxZR4s05b4r03EkjV9ZuOF4ZxjWR9pv4GSYe24zE3eS73BqJh8SzO10ttvbP+Y1X
baheMAdEHg8ceGzztINbU84ZaoxYteVFaxfSJHuFB1UWODEIEfAK/LNrgjkAA28o
smFUcVhK8+wJtEDXhPjLvQ3lA2HdaUAM/atcqNgApLGDze+MtminQP4JM+3nfP12
WkkiwLf80kD9wzgj7xs42MbgCgQmzvZZtX1ZlzUoGJ6Jsp/JNq0rLm+mGQaV1GvD
CnuAMRlDrIOBt/EKO6QcfI5tSGvhVm00cz9aQcnCn1b0dQ94DXujBjurLi9g0dvh
L2YFKesWZoLHsm58CFYfCFdeJXZZxd/OAY4W9lMxrcfFAJUZATVfEFsJbSTCbPAN
pdMOwOJ9Y+apm44p+d1MEj0kZMgirTto2RtxIOZlzYB+NgLekHktFTMbrwL6V2fS
XOSxJbLhSwLFUJJ563Y9KBhj0F0oJhlip/GRRGsQKFTmGdX4UExQegERQeu9ZINT
mmzJxNECgQbOs/Eez+Tykd7IVMmdAjyhepOUgCK7ZppJ1ch8uKsA8BNO04zckyh6
B5LH4UpZAn+iud0RWVkxbO7u17Nljeq6wQkQovPMbApeu4YsTvNY0buDPSTKv8Sk
WCUKNUzi2cSsLeS8OXBuNym12NHxUAAVEdI2+wAnrIVEylHF/itOSBD7u6hV+JpN
evKGnzCnHLzlVU0gNURlIqacEUxdN0eA5JAqAax2e+lYYpJRnJnIwuxLspGK2v8r
U4xFeZSsUoCewVo6IL6yYHprddurKKN5TJNQ5Z0d3o1Uos3vl3e7hjj8WxvvGgnN
tqrMyZ4trRj6GxFe3UGPnWcnWd7RNg/bqA0k9i/KeLwhWy4PDaIlFc7G1OZ2nn4v
0Nj9th/wbaAxt/N+k+nJ9aYf14weZkHNwy0nnA+qQmibduyCw+dgb5fxfHAC6s0X
RWkm7hhJKzi3x0HDmxBQbWJ9AuSHLBBGWHaVRqu8B9WI4pPnrnvUKypy/dc/S5sj
emwK8Gn1BTdj4l6bzJRKD4hyXtvzyRtnw52Io5hMhI/1v9B6uLJ7TJKIq7e9eW2S
61erxDnaAQd8Z+f0uyQRNJHHhgiTZape2wzkeO+xfgiDB3ilQKtITw1HuQTdesWM
qR8T1vVZwLAdM5unpdQ3KZW341QUex2ly6Ipy5aD5lZD9zliowsaG6njT/Jt97eN
ppjG+5h+rkekIxNMt47FA4G/kPRUw/7kz2LJNzGx7vNisro8ccCi46+zvLYqKYYY
vefQ9znNt6+pMbgnE0blhObSXpD8MOvvpepUAgDP+xk65PPtoLSTjNgG2CT5Nrx/
uOe/QG3To2Q4ieTLdvbz1bB54/8hp0Tu58fz9eG6AVQp16hhYI5nvvZBrT5SfZRR
Ud1Od1LWw0cuueOfIAzljgjeot3fF2LquLzPDg+n1dW53ISgLPD+AIfVFDUVELRs
UAgPvRI4xg/2+W+fRfW0wuchjRFtDIvazmXlfil/AEkFxgewXc9eM74dKc1mb8YE
cr3SJyGc/t7d+5TybiKJ/nj4xqUf/LtCHNwKl7EOq1RNmXQ66OQsw5URohezLTy2
bzu0qb1MdDWaz+X4/5ZabfC+RZhkt0jjKq+NAgpXx7Azxf4lypupm7Qg9i4kbvKo
IzdBlwIOqj4Tx8wvynbBmFYkYdMVISsRdHnUGT4zOB5G8WjqgW7jvqH90N2VPfGO
/YCpr2Nit5ArKF+6yok93XXIvQyk0cM06kW6mHubIH5Aa06d0c7dSX7ITJFW46G3
/leO/1EK6Yi9o69ltN8yyoGkFU/1MpcsL00lnz2RSpuLzX3Ltkm3PoE7ZHTTsR1/
0Mm4m9+yvAQUxymVOOz6Z+/wam0CqhTxi9TPQ2ZEK4GHY4sbbH4zCNMmZwjl/l3B
4UAVSt2Q0O9qUJkoppMjRqzTpQmRilbjG7qMMyh0TIbGseTGZESLp6/hEEz/z04N
rCgNJti8tkiSHcNVqTmczzdc8R99jU0Qx6WgdIlk3wRIMMrocff++mwX71hI5fCj
IUGpkMA3vyb0jQk+6iFL7wm6Ub+DwKmbzoV6TfwYOY5AW2hMNTgrR6czD8HHccDM
s00xzqI7MYS1wOYrFuaEqW0G93dnFp1Gd8bxVfbt7poYjzdjqYxNqYTE6DBzx/06
2DX3lMTms5xqhBPkhDisnx8GyAWsKRiHJuzw2GVxSjC7Vwyp1rAaRmSISy2GNGbb
G3htXXDAgfJ19TwXZJyYWju0Hu8a3oYajI1h7MjXQ7mKLt+XdAfjFjvQDgFL3Yk3
l47wu0wgKiHuvdKylAFy7QTYQ3QqAZWRYvFF4XPmekfgQ2mBPCUJR8qcCCfxR50v
7U7w4LfrohkO97SWPHY8HrdcOth1vQRN8gWVFQcXs1o/NvX7hWmGlR8njLKRZyUj
apbO/z+xniQ95qTpVRCGHng8zrbNEhcLnr95WQ3l+pU+tAp34H0IhgFwW9bgCqgD
fIOo0AyDVCcSBa5TyyYsxpAX+HwMBEogNlORtmXnJEt+MhWAn9t669zP8RNNhB9D
Bipq0dJ2/5BseZkaDUgMtjAVFiOEZ1tiYtxycu1uyXou5nC04z8TI66uP0X/NGEz
oSV1cN8iKSgHE6WMc22JFjcN3uDbg2mVHLGF9K4JwdGkSh3xKTmSbOfu3Rqd4QH+
ha0yrDszZ88YJUBEIgGwiAYzaBpNem4bSooeHT7KIGxsm6lC0Ez4sLv9kRdtQq0L
O6AfDpko8WYLAIS/3n7PA8/dBcPflRrpPtn42vjcBo+dL3YbOnPxI2M1OBfwuzI+
avplfrqfB+B8vOWnq4deMieF7j5eih2JeXBxOxyHQTckjkKMkdRahcp5j88UGfcR
x72vRRs2MmUlLY1O9uKeBbhDLDdQ51OJb8iOy8yOPBP5KHaJVfizOc2auawTmF0d
at8orpCOBir6HwxWEZXMLsAfMLPgvsaZqK2TUKGYelikcteKh8pbJMvLkcqvrCwZ
dXbA5GBBWdpw1dT86erjdMbs0464l85kCrEkIF7MLyecOHzqz387tyF3dXpItcHC
5+LVK43A6gUTDCSUjQ221DjM0AALo6yuFJHApKkk9GnJ4il+Zj5dFSutxnqF9OS5
5iXUGhw+2d9B63F1wb23Lda2lsOyZ6UY04lNZKl3523Tzb2zp3oan0M2gZvexbjq
1Lg8C0Qhzr0VnAbUgCjDdlwqK4M3cJj75GwPgPjhoU2wI3hxyA03j0icfeVvXghY
fIrY0YLZ7X7m86WedtLGOqUqkurMWU4DQKWGo/dB8cAT48EYi5HWqHDLHMMwDdIO
JJ9j4ZEKWS0/86iIo1rhssfb2od6uqWpBa5cSB19dTGWSoq1BqzxuSa1T3Sl2oFZ
GPdCXBnKPAaSlNHS5SY9OQ4EYxBdzKxMVxcXsgb4oXDpwiND0ycYtseTZliX/Xon
RusYsmDm/vP7Ff9wr0dqrkkubbpzVfGM6cMIJJ8f7uKe7WEz99cLuZcG2glK1A1k
0t4sn7WCzJwDUmJKAmiqTjV3dVxkLAv0tiOxeNxpUiiPn1bJP22t+DHezIT0BM0z
hC1Mt36oMh9gKlI+Dn9WA5aRNTbFL6Vi4bTCIpTzW0UCKmd5PZpAJtNTb+Ce+mGP
vNeiquCP3ozOd4xNEk8GbfEQc3ahNX7GzBR/PkslXx+ZwVYj2zNs0oTDNsIFKJnM
4a564ZCFvKsh4IPYqLyTsV7UqCDFk7IJik2JF5zeDlqM41m0TWQVzj3aDgUdfN0H
Thr++NqPBKop7+ithVYsPMHU2PwpvjdK/iezr2PLhSlRbDGeRh8UCbBah7jsjEvn
zYqXRdN4tjSW8hkcJltRAJV6ltXPK358W00pBvOgAIAX5j9UnLYHMRrUDFiCe+Hq
VLo9ZVWfGr4tDHPYu8vTOp2nOuCGbAhLqOEIPK4hBqtf1P0pm/xD5WnJmy+o/wBh
shGODoh1A7PcCDNkt49ObhYuAA/VEIUM81T3n6BO5rtkFVEPV7OSZmTFJnAisDA4
B2Alz/Cao6wW3ZRxUE1Y7ptpYF+YNklyQAsT9ap8eBsXwuMLW7adXK8QC87geoEY
Qa3bqmjTpulyRtU6429kMFGSUuRwjZ0Ktt8uELiwwf2nRFFahIShIRpeNmQOoCvD
ysB7HtJW+SzrtdbPQQ8r/PcUdeohvwPojibCoBHirRrEAyRBaZ0ccVnSfH1EBLdr
JHQrr1E3IRw9y06YEzglN6DHyyDeMb6e9ikcT+Ye6e7A1AzTS5RNh1qXSQZs0iZS
lVEYcvSjHWUA1tUXuIwlMeXCCvTRu5nBGVeECiUVQKpHa0wh+vE2L3IVDluz4AUo
ZqoYZ9Jpnwgz3iN+EyIfx8o4k++XxyVJTWnhjeigLy9cbgEAXcaQERyK8o09rQ7y
Cu64aq/tO7Zssd2dIVoq8fZSIkzdXp8yTrJ6zNOmsFPNeM4RD2kmwZ2PMbemTAAx
Lpm1N390AqOPtCWQJkIZ5D0TakVi0AYzKEFDzWp3XR3mhuTI/uXfM4m0oyjD9Ii4
/pPz8W+iqLx7Y0EfSfSDRuMrcbIXMAvG9sFOmkKCIVBGRufQCthoFeqCgiJALBja
d5vWaQilpX9ESiXsBK2G+JwgOC0WVXp8lLRrrMFqffkvFlnZ5KFegkedEkTrsdxs
HdAJjogmksjWG/tpjlQGQ0a9KMnlWoWlthruOEAAsmWOk57hSZnAW3SECZU0r8Hw
uJmKGHTtG5HxrXq0yQBSINV2T00iA4kDKfUj7SwnuLTuw3XEYhECLc1SI4ytHww0
6Y1ODycWL1B8bpnMxQ3BCrWgB98vY+NSTwRiGAK/PXL/J4mSRMPOCcHR5ye1clo2
z0JiIYoPASphSP+7TL5T/nztDvUmpRYs5pSwdjOHUjsaHKctZyD2XBlQlQgWeHyd
Otvcumut9KRzg5kSocmIl746ikP0SmosfNCvbmzYvRsRc/HkcBbM9iT/TiMuPpNj
AkJb+fRdjWSEq3EeKfdlVGsQ9bbal3QmAHdgUPrcKXSKO7vo8bw9nN9WR+Y2Qcnd
UPca1X19aFHhKjkHflrhPAgDA2Argpg7C+oeIivPBFiiTF9tot0ze9aMMvolZjsQ
Mkq7wWqNtrGzE4po7M+1CbTmhFsNFQFneOMp8HKzmk3lK9+llx0S+ThbGHhc5biD
k1vaX1NCJfTuG34WvR//GqWGuSOk+Aq+lg8nFlrtIOcOHR+7s/50jwctVxnSK+42
4X7o5XDmE9gQDeeZLISeDzdiPfo6jeakvSHy1ZhL00l7lICx94YiNB3tBdLDTrkU
T+YSO/Wz5R9dDrAk6ezUzxAQLg6HInsoQql/umov9XPEwc6gamODGH8wm8Qo8zJU
To+tEnpsVNcYjS2bnma45JLNFBdN06smuh3Z2dkthLkv365eFTK87LBK1uPtaee5
6S6YDsKPtzY9vqUClHwl70dBYGlX9M4IirZNi5qeX4XcDZ8GvuvmjTf8AoBOa0Er
8UxtWWrFe0758Nprra62Bs3XWkJw3LFxe2DPezEUoq0QnPeuqPfDVd3CKZjV6Dmx
Jh7E5eaoEq21QuPpn1565zSut8fSEp/x0UX7ATeEp/oADHt6baVBblZmBk5tJJd5
248oeiULPMmK5ehblKWziryUvyRHIkPd31L4odPEnkvczFhpAfVj9sNQGpz+in84
Saum4Mk4aihFMbI5Nz+1MU6isotv3jGc8lVWPn5fdgklTJp5efNyUFyYtJZiFqdk
7s4DTgEYndSjyNrJBaZniswTQUHV7M28i9HzW3MFeCWgGlXoeaCq+8WkoRz/6zUl
UMkMU1JXzaxy0soCtZHQSU79Va9LACZyrN72Yb6PUWrErIgmGsEvHKtcvO0x1643
eSqTTD0/B8HgIxG6Ksq1JZrj0X2tmkixomiTG4td4iSX+C78Au7U7ncUdkNMAuip
VR0Qh9+jNSqb/m8wKX3BovMyEH+6FH3Ff75MpqLdaSZjpEhRvXdPkln5ZTHHRNjE
LZTk4N0emCvI1JAx1zXQHDNadq9TFbevLucOsBKzDSVkY72f2G9ay4JBTkqGn7n+
xr5Oz5UrUlTyiHuMyYfDX/KS/empnBN4vyGKlRwSx2Gdqr1805rh3M7U/espUIWv
/jlMl2wGPkVLH86u/wWBwTg/IL1YZT+V1iQwHKAT0v2U/3fWxTzZjxJf3l2DpzyX
5V44EzsCL0x/Oo/y/C00RLy9AcpvEHJGz1pKYl4tN4FQXkJ9UcyJGHLSgDDD4L85
/BwsQgJMYtkxioufXtIpyDuVdNjqEejKqUusa4m4RoxLsM7gkqIlSkYnJyc/FLD7
wYKktQwtX+abJU9QcwiQeEbRXFMLcVpO/ds2UYxLw8DEYPVCfp7nHD5ROUgMCivi
Bn79uSO4B2nLAJW94byAhmjqUbzlM+0tpx3wS7Et0y3sRR3cX43W/plXQiZlG4yO
9JwokW3AwscyUyXKV/FwMgXsZeHzucRfzQzSkuJPqf12/xIHcxG4VQgnFIkb3fhU
4xdTwmCAS8IR7kV1EXvC6DC8kK5TVX5kNeGkM8gkzXONqB55XteHcOsE2V9UdCOp
C9Z/COUn2nS2OLB8ZFVnXqzDcuH+CFJEjokW/2ZjyP18ppIFoBF8WMX2uWwgMz5V
MJgvOlYcHxModXeuDTETVEwfH7snS9qTh7cTlVFGagDIzX1BE6fRcgplHHfdBRlB
rnr+iX0XmjyRtnADyF6eXaqLRSj4F/HwfrwHreQ2m50glWGLY/7b1dcm5fz7wgy3
BDDuAl2hGQYOva+XXzQ/Y3T8N7ca39pL29wYvnr8m8tV7kbvo99sUfYlhGaCmaxj
YGBgHhtEnQISClMOhg+/ljcc72A+uV544QcRIM97JMK/2h4zpYEOx9yTo3SJCK54
SwLKD6o10yXPutvGk2ZtK3+yiksao+dRpfrAFCwwOqsmLKYDdemI5IOSCAa11LPv
8E2Ge5aoVGZfDTtdAhGoDOuAQcVxZDvVKVdB0SFgXl3daJem+6INqLvwM8tHH+Hz
sgE5brJOksNWNoKn3pzbvUf6dIdOS+UNF6zE/WNdYkm+coSKHxLV0SkaGtG5pq+N
yqXUBOxOPSnTbm4ZzBZ4Xr3sWi1k/TdxI9kbWemNVTRfPwRAHz00oiFP3H8ufsIS
Xy71bBk43MBtMYZHKdcylxnaEOJnF5eFMNEB8KXftdIEgvuAVwM0d+Nub7JoEXRj
7TwOetbNfgC/G6R7u5ODknen9LuP6/lbJ5HF33ZF6XSfKXMrT88wztd7VZyDs/KY
6qXWm8U/+H6C0oVau/6jP5HloJ+uTZ5vPdgBDmJGnzm1XEOCTjN0Lti6kZmolHTV
nSN2KKNAAlHpnW0Bq8NtR/J9ZVhuLd3ZoVpQPs7pT5ekFot6CKnenAx2iV6MD/NR
G4taySUV+h6u3/721Pi8FoES/zu9lQh2WspmJX1c34hltxrdHw1OwrJYzQVHVhLy
PI+Nkv3+QbuTVyc6ehxVXcVz+K4bQXeD6WfinYdEqd6CIljdrXO9Ek8LKhCz1aJ+
uBWIx7fPnyAMzTJ/UFdCVg5mF+pVcu863+uNJXmkSU2xKwK8DIm33CTm7kKwMSW7
Fg28sxLIjTUTS/FvkOdwGG+Es7xqXyRKIVazv0ndZ1k9K2Lj47Xn/PrOudqYrwW0
22PT9xGg8urV1ZFlB0KLikV1T5XqCPlBeze75CYinyyz5jGas9TetaDZcz/CdWJc
bPP8tNz+XW2uTrQc6DavVOsIzkw2lxJ42tUBEWNDzdZiJfPFnfpbujU5sJaXmAYT
ucR0Z78i6+PjbSfK/60FKYuw1dVztyymHroLHZhZcXB/dBWjP9eevxjelW62IXCl
JPh1PB2bH6WrWP1jJHT5vNc1zywueYcI4BG+qCZvm3jy88XAovUWBSaw9Dcewelv
JDNtH/sJ7MPK3AUyqlBbzUMPb3IY7l64mNxxPpnxPNJD8K5xfd0fdbFBwbuv0hFJ
Mfoc7bNcXf/jVpv0G5tAnM1ZoulGI5zlKS+SgUwDIT5lAPtMjtS2hkZQrsgtGACL
HREtuaMCTj9exyCMrHlZUm5kJaNTvj+FVwTGiYZIKVBEGsodyyjvBmfH97CSjJEq
4GQprA9zP7shoWDTmQK+zTCtyW59J7DEWPZkf1PKY/5C37IpPbgJ3GzULloxI4Ox
byewzA0utM6VFSTxXCsrWWcnL8fyNJN6zCJfvQxUhWPwg5h+SDTXum7bgnFCMozb
/6WWkKMD5ivfTiBh2HTnF9uXFdY+vltaVn9KPmZBKepJKCV3KuimLlDhlR8pDW8j
pQ1O6HujMpGMLufXfoRFcb1S/9tojxKJ0Eu8HAjUUFje1tcdRSRzqkiYdPCq2a3e
G9BfzAWIvvq0/w3ZuTLLdyhVaDWK8jNXM/sJw491HgJ+sSYsUFsrpF/4WIwvy1vb
0+EdNyQK2gc7ggDWcK+hDcJ9OJfIlGvSF9B3E+nTtei8Rd39VoWquPC4F6MtBz65
7pc0JFmhNkX6sVUfxncy461anJc+DgVzP9j7D3ctN21tc0DFKmnHX/pCdgmPQqB1
cQKMkyxYgFH5QK5vqd/E+eR7b3Nj3FY2FNi4W7ss0TbGCT/4jWP32IntaquXm7EX
mDMpc5eWeUKgBFqU7Vn5vQCANqkVf751XiZDC/agpTZe7QOOTEX6jDnDTwIUJLj4
21ssSSaWl4OwwUDDgOvm+1R9whKq3SNSgXA0MNUDIR7csrck142efQ5dRWY4lf6L
C+9Yw0WYm6d8VdaWun+RqyYBczq7F/H5I/HoCog0mon8U3eh6r+CfuJnbGjrFjYK
oujmtxljJI+RGY3R2M+McrhyutOEtF7YmypMnRQo2sy5NYDZeFhFYl73sK7nPKN9
hMq7vl1T5ZJZ/LLJXpHTy+arPlgzwaskxCRWF0tnBNt877glFBOX92MPIgEzzAla
vJxf2YQDaKLGV2NX0Yyj3w/9LlUDMsroLuGYckcOKvbUb2Le8Ccba7ry6DQvI88M
VyAdLiC/DKQWgMABeCWPP9esuPU2EWRn6fuTIT5/usgGNv+oJDoFEJEbwPMOe0si
F/heXJxVOai7xyjZu5c5ULzCftAHUQh74KK43RRT/x9JIUhQcaO4IEGBiXl6gB8c
s0buVP8epjR9NuCuPeO33wLGFKDpf5n3Ga8EI5+zBpyCVCqbzhqe9sS86R27nM4e
/rUwehr4h5pVC4TGi9NZ93dAW/ibrw3fsgCYaIKOHw787yOiraFV/Z/MoFMfAUNM
pmHwHIJzBxSdhxyGfdGc1MF28AzanFdejs+Ef01PCYufPQ5SMIG9eCyjwXmViw7Y
LAcA3vZgY3/Q8MBzJVpXc1waLlF5ACPZQxr58UktZfMVnASRuwTEgnEhNgLl4wa5
zwcmnObntT/Gzztc9s9nllIeiaQLZAaHOJYdSYu4PuMbcPXo9tGTC2wJsfT/eeK4
eehCIH1xsCAL/HNpcT2o+Zi+LJpX9GIDwI34wV1Eh+ZS8ciJUk/4XyBVS1WVqRP3
l+MSH0YkCWsnI05tLTJmOreLsNaUgxbVf9Vj0gLTFFt2jzCUZNNnLXm6D3qx8QvA
wHL5a6bdIg8FD6c8eC5I1d8a7SIvU6iWoMcM7GGEgTwPN9BWVLEOyMt1WHPXK3fg
Zat8B2b6zp2c3W4GI/6gpQ66HUAdtE9h12pFzdEGEUqN0jPbwd+pyWwHodIW/QlL
iS3usp6jO8ACvddVqB2uZ6vMV6VVJ+eWQEQWwfaTow9s7i/Mjm92d57jPxf6DnJ8
wCnW9hzICrXFhbJ2tBt9C7sv7P0tPozvzYUELj5vm0DZI94/HdPmqUomdmqFPMtT
7GEe1l719rKQMMH/teTXk+ePE1VXx7gPBzg36aLxPYhzNyWjexyKydXd7zDYSK8I
CmrBQgcQFdzVyAKjO44AL67ltNy8GKjAiqKSZ8y2Q9S0AqXcsl1F3QKCJiYD5tBY
uZ3eiG/XTcULjy8hxrJ6WGt8TYg4AY5/Qa+gcIE0NT62HpLUfOWfAo1IEKmiweta
PxK2HcNXzscmG/Ccu0xxA1zSw4ICw+i9Dw0ztSWp5H+sDWijaJVONvpDAWz2fFz8
tkP3QEf6qr3smsO1IUR7T2CnGaMDZ2FQXNu74g4tp2PTWnhgxp8f/Kqdb5AvVRu8
JuPzkkSu3gJIJHYQ4PDPejP4ltXFsmslUNFSltaZue/90wDNNcifpw9ivBKb8yK6
OiSZ+DhPebXnBlESHZ4qgKCvbCZanw3vSznjKezTPY0ND95XLrOKYC5ckPvUp1G6
MTiv+wMONrRR5DjuGl6AyjNAS3RVn1+RupRhVj9RWrNr1BA0Rtt54ZiivtuFnyyu
CfPjaQXRjq0syzP8Ik3p25EzMmVMHE7vvVKvbGXvQYZ9R8u23kpLoi0wPODV/7cO
YBltnf+Amn1zcY0ptcan5jl05esoz1gBhdSHjiHT4+rixPBZ7dEGcCms6eyeaQc1
tCAkvyPgrig169TozAXNE34fQtg11AE6l/5C0+gTRhqIVx0QggC5wJXKhZVaNayh
FU1Scv8bFOV7qEtDYjwAyweEaMcyiPc+vCgkVQycXgTIGJHJeME05FAY6ndd7MpD
xbsPnch2IlHkJQaB+kRzcSNGivqECIwG5Z8/F4EfV62XlP7CsQXqRUKKo0s3hqla
uD45qDmwaI/uLwSnS3Z9C5bAxphW3nCRiHgKu7ERCddfu+sq8A37EM43RBSe/lZ0
gwNzepaRajxu7HlrQ4KwmESRpYXAtcUistVg1q5ahGF8Yk20MleRQm2KUW4T3Lk9
uu5at4jHAIgW0ZPkV5w6Zs2dZ6lEAt6QwEP/6mEygydCy4IxWd3jmOKo3hOLnIFU
gZ7IDk1pqofs1e2UYS6zjU+xMaUvvEzQd7gf9NkAK8LmViWMu6n+p62S8h14Q7iP
4N9FiSBZ+OzIbbSIDWzuKmaPBrZ0syHL/SzxG42IsFyjXnqDgQoCh4PETWHCkOSR
tEP+fmCnazoy9/UWXT87kkG2Gt0cpINCANmjJ9f1AghcV/ozKaANANkch5fvNa0+
X56L/GKl+4Z1efyLRGuEzb+eqtz4jTM66jMbwwYrwsrtIeQmFIAJ7NtIq29e1hxY
ERHufcE2cd8xBHcAkJhrYJz38whZkra+xq4T8Wnv5O1yPfJjF4lnC5sxDEQ8jPW2
LNEH44j84Y+kFaGVoz84Pb2NcC2gaBBL5TxfjLGwkimrgIErqVTtrx1HBeYMI4lV
jnhgLDzf+Ul28DfAA0czNrrGAPQjCR6N3ckTk4QTNm1/0eDXgsr3qWvEszhQHZJ+
Iua7yRwBs4djj0mMSv6Kkd6ydQp+WvcEdNDFR2pjpAvQg1+p6m0gi4miHiX2sOlt
Ho6HckKsa0dKKuCoZANbCP85VQMb50pQE5qw67DXcaJVg4RPuYU1+mijmbrmveHp
PMXcwWByIbhrbKt5TpE9OXDIVC1Z2smxwgh3dmS2tybWB/z8bg/qsqqy93pdREgU
3TMF0DeoNfMcLQWBYQAWx+culDfNi5Q+OzhLN7X1L37rK6JiTiz4+C859woTq1p6
qwPgi7a/Rqryq7rbAt98HaqaBTItI80to7krrFlVROTGqhfWrBGnMSDnwWyLcpRb
u29p0jd9oiAN64uFSrJmUQrJu1YCd9w1/DpF8Qj6ZE/kkz+CJfrtjKL8Ij8xhUUI
0DdeeoAyxjM6hLp+VS1EO5ClRyg48T38OiBAjzAsGIOp3DC7S/g8sKQonjklocWG
i8+pephG3D3BAApbYx7khKSA6KVr5MmXkf+SHeVHAzYndlxaTTpIGNMjC4BuDb8/
NDleIqCEtvih8IVv6DCOF3tajh/WSgsGnLrvyk/NN198Pha9ZvYGH7SRIBp3Ki+J
lci0lS8B+1IOFUk8cAgBTglCiGnb2YWnEUIDRebgZjRlSaeIOLq/pcj4dmvdsEGd
t9xprX5SXz07VYMmbv6+lXrswm3tm6ry8cm5HWNCOMLpitRBszYP/Hz/msjviZq6
omKD5VB0JyC6gHukrdHsfQghiuqnuLIS1ZXU1qKWy73GFsv3vZgY7P+PT/37EBY8
fjFuGewVmHUoIlxt/vdmclE++Gc+mAN+iY8g6VDqz3zx2OcYYHgKXHaVd4ZkcEMC
ERBilSABXTfEzn8grETGIwT+ZO9fL9drtdtPmZCVHGZpN+lHSecgMs/nr8rQr1M1
iT84CBBPp+Xx5DB19gaS8FGBJ5W96IFQNu/JHUPEgsjdU+EIqOJhiEMaSSNIugBt
9VzZklpQYnRSejOi1aLKyA4HS7G/SdmKL1wYBrcteghtmyrnx1jeTV7EBwwqIZGe
+O0q2bUkQL1RMwAmWeK5zPZyyJagbWEGALGdBjXkq+K0flUUbUcXl+ygI9Mg8nv6
tW0zIz5MtpwedC+pagQE5EWq1SGbKvWrhRIpDoH3vTkV2AzkscqnwLLUfatjECCz
moCGMGg8jvaA7sW/yX+zmUv1SJXLUpgu9jVuQi48DVIqgxtSQu82HeCO8P1id1Ow
yAXVf9/oEes6vhFZXYMzDzAEprojv9AWz0WFzqIdyDExfcNZzeTlbIwcMCUnoiA9
JDwshhajBZQrJj1dOym5ZGEuSpU/dok8ezeCl0XMqiNJUhe1niIguLqn5LrK7haG
XFiyQ+WSDwahGOz1VpM9bb+QnB/iGKdbAkQz9wqdfscbjHH0xGmr9l9gyNNygKq3
x5+kA8bGJ2d78LUliy0crJJxzqY6gyD646M7PCRJRxR99EcbFyA0DS1KN/aIS3uV
Tydgbd88iYz23pe6LEPz474gTeF+QMQSu4uvotxmnWUKeTJFZMQ8IFhfgcjuPSLf
8CFu9+UcKDdAZfKGRdHTqnPp8wEnCWdIyqXRJ2AgfxthNTgrjppyzrSJ13C7iMv1
guLnhAm2Uj04h4oXVblcc6SNRfeGK77HM4nm6HiLPPcXurUU2vLN31mua7TFI+1Q
1LKCgaUxNNGcoigXEXGTnZvL5cs1NBFoOCLCFdRJKBsyqtLMXhlpUFmGrdZH00Em
fBcdgd21FqBxN/Y9i64P2g2P1DNGWWUJ1kbbd3AuLSJUWTb45P7yCp2V6Exh6Xt5
XErC2E/6Feo6VBk3VVpn7qBSnQ+lKHZ9n2sGA3ocn3JKed+ULhvGdtGJHMzapwWR
goYd8+0Iai11D2zd9hbL0uYb+w1dr6IdZz1P5DT97CFN3mFdUjYfMC8yYzIKM6AA
+kXj2XcCNX1QJlxuG+v50dhxWdldARnM9lXWEoY3V/ihaai7c2WbqhS4kF8XS0jY
yesabes7pWrwjy0aZQMt6aEaP7gdCGLaqnWySzJpYeZ3D7wfl/6GXzaJkUBGX59N
VIoWllpXmH4KSCD1NVNN/lsHusIO13Ul433HiIsSDZGadpQsvsW3GTxTpsQJ+KzN
9HHfScSeMbdyBTcugZKikdxKYh7F7PKbwe5wzMt2gbGEVDYMTyrBnU4d6xUUydp7
CzvpvFnAZbbC2XhryxbnNv8gDjy63fq5Do7oCZK9EvSeNsubDt1Fu3euZqn073Q+
zeSlByUyz3m1uI8LloT3RzPtpjMekK1MyH/wGaKSOCt+ACQ/yrrwRideEmAcaO29
qVL9XL6WbFN54Y3LlsEPW05fhuxymF39Q7jfaZtCDJajuO7PY5gehU9eomM6xg+r
fYwZl3DeDCtzlqYoG2oSPjrEHT+Qci5+RST6HIschuapQrsroZTYRld0MYJqslt4
a18rTP16yeUK7TPsfqj8Dgx4PgVkSVXbJSlbnWs8k3CBWw9QOB7yi11MVfU9bSos
KLRTQUDycsl5PFzl1c5gX5uy3S4NCtaJaJNHxVtQeyJAuRrDd1nnGf1RauPmtkWX
lXIDvztU+Z3ymatzWNfgBgmYXOjUpYtWuN7zy/B8YbEtqcZXJUsrueaWGV9yOpP/
YPgJCRsPZfTek85NVMq6JAopxKcX53PinzailskpgsAxk7pW+n/ZmTJVU12sqvyu
dR3BoOLKTm5ikL4Hevt7ygxA7Sv12W7zpDdWx5WuP1oAirLX8D63G5dHVUfU0Awe
LQSj2Qj/IH8rbcHGhohudJpPXRvgUgb2V8iv0ctjvy/Xo5zBSv9XEwHJcC1Mf4WX
cCP0SpDl16vHq6BsjX0MZ2rOtb3wrwz1ybRWYw3u9VMsar/D2m9IvMbttXFWkeag
F3wdOI3M/3woallNdOLQI/eU2NCuHQfJ/MnxGFH9HbpqFbYJJVPTHFErtc7h69OX
Qr01t/Moj0AqXUeEvRuLiYkaJ3QCtOHw5DP4eXfZmFi8uVYHIjtUka54hrVelo1o
UqcF21ohzr2FZ/VlF1PYOey0GJN87KzElNA6GcJgJ+rTLz4BSa86NDmHhDVnSl6e
DrxW+K8ykDWlkZw9TlcfbKgX0Kf+6xgcsFEXYIOUgH1VUYhWpFjuw7LnHqY7Le20
n6a1on1GfbpNQ5kofMT/gC5Gj0B1n8Hw4ud+cGxS98FC8F8j1FM2BvAyBRPSPPYV
2eM4t8j0nWt12qB5wuoL5WcxNuGr+Lqgv4I+FYCvlL19t0odozDmPn1mWmYFL/gQ
GVct/TgH00/VVOACyBm5YIoGEh868UaMtVTaUsz8/5dICqfaX6iPZq3ELiKOrd3J
I3exPFBRAG3CqesHQ0EqA04BlUjpllI+wwnZy21IbHFRhKC6z+UDLV3KN+QamX9V
NBnTa3cOnols9S2xCWIL1CG+gx6ycEO1Gdh/t6Omc02FHHSBnFSG16qwmUVIL+2C
VQ8c6W2xb2qSdQa0Rz2bZK6hnFkhJOmhLgomTiVT/dAAttwu81sIOKmVorXRvCsa
ApgeXYB+FlXKmbHRK/KS4S7QCAshqUZ4Jo5aTAGOj2obSkimotd6o7R1o2dv0pN1
DZ5+hLfLeupY90ioXiLifjAza4YKf6t2vFpTf0poturuwXfi8FZa6TMmh15r29tm
8rX2WdD4VdYW86daFqvs4VUCDXM2mBs6j/ULA7x8L95lrsOid+Nznkb/Pjg3Xx/o
juVMCT0q3ExP0MHjbS7e67Lxg4eV9HeF8k2IW8nHQZiQKfPlei42u7OaPTq+4hPq
sHODjXs1Jck5D6I6JnrF0+gTxjYkB4/LVTuq00jBwy6euowAS5nJvFU98/LrtxRJ
mv6Ekj2DmLCWe0nvPplcrNa3LqyA4orAyOQ/Lq/o/+O0v9U3Fj0jBl9tjz+vFIZu
O38GQIq+HQJP+4btuW+2bq75wFrxszUZfnCN8af7q441FrfAJAudKiozWTuOgmLV
8TGUb9YJwRw9x/XST9dhWy4xqaTzwraH4XxQM/nfnRee/RihiWYHxEni8hNtH5ZW
Xq9c7ymo3Akx/QJF+jZeDQVEr/u91gBskhPzZMBYKsuNhq6IYpeObZmtFMgYAcOV
ReVQH4bxlW/i/WBfM5gFp/9+Z4+DT/OMXWUVWjkhgG8kDCzVW9LT1bXQpp4o4/56
8DyWusXfhHPrIU6A3PVkCs/ubzWb4hioyFGVH1XXaF+8UcnuZlxqBgGhJwPuRnWv
hO8rC5L3s0qkpDXs+g1wncRxXwqoCzF4b+JBfarJc2ZaMxKTsr/JecohpfagF4Z7
8uk6Q/fnZwoMycXivqfMjK3KQSQ4VfywFXH7qDO52/iT0WftS5uizFgauC0Cyh9l
iJ7+LPZUDTprp+e7HBOxpuS8DCHjGyxd6ACiaorflY3T4prTV3isT2rqxkccJtln
S01n1q9g833o48bFWPYNYvIJsFV1RPNACTzKdtkvY5/Az+8c6mhKw3EZww9/MMf+
w2DDkTJieUl2235TxzNuIID3Yn9OSXtbbAH+cNwRv8EV+s8Bda10mrYeVf8qqHGw
ZATslcjtysIyxaYtIoqjshnJnyjdfNYG70OIDSSpCHV/EXruq3RKMmfdgDYi87rH
+o7lSnsCtR5k6Uxop/9Ouiwm1XEtU0aGCP3p53ytSDg50WyIK4TWt6wPZiGYEQ6Q
vsrwkAdr/jfrZRhMEt45gSjAi7aglMD1kPh18AqqiD8vOgzDpjkhpZ0xpAT4dFvx
XO110Z3ptZ7Zd6u1G67X04dmDyQ9jXaFOoa7uUFNOKdlIJMFmmKrbfH/9p3zTTGL
Ylxsw2RaFEnlBP4G/sA8/H75DWzaNtfzGYQyt2gYr/2wjpwME/L2rAtWthhsq5oF
+0nDRKUxgOYHrs3fh4wnwGd3BscYi4A2L+I34b1bkbP27fxMKLgA72/D6m3TOgdh
EL2pNzgk6cth3fBMl255q1iKxRTZcx0ifpZEtIBibf+sKRc0/g7LQObgvX79KSa4
xwmhf1xOoqwK2FoP9HTVJE+T0WlkzjBFpvGbentnUpHpBebSU5ypswg6oELYbpLn
XKI3jay+4bPZklccbhorRnS+b3XC13YYeg1cnEAKoPzREbZ915Ea+v/+Gbx9ON19
/20WSc1NiVnuuvnZLTd1ZbJjXzAt7sKEM0gITuZgzvrf+psoCFGAP6RclEZh85Gu
X9sQ5Sk50y3HoPafqgI+a6CN9xHt58dzxfbqpIap/y/DT6XbdYHuvqiGQtFzny03
7V4ZYTQDD7hetubh/CdHJFC9jJsrkXx9d38LcCpzW9X7K8sD1Vwa3sQ0mUvcTzJM
HlZiw2+NqPFDioOe8nq8bVfKTJ0n0olzG+PGBpdgMpmVkPhXEa/kvA8JsfkSTgfs
lnOENnUo/6NCner3DOztWatUsUigTehvN1OoZXP1WX60CTzCa/wX42HijN8YxYaD
7OYaocnOOxYHF72ZactuTdgub6rLMLokklBgm+GgKsfxuck+CKizCW0ZPJiR09wo
1EFfZEweHncFg5hSfTuKZsI6awTTkSI1C6GBalHx4LEVBh/BKunj+Kyq/CdhxpjA
/4wYQ4XqXWQE99eLoN0oJzV+yQeI2mKXrPUdKLan95T4Fmaxi18ziSmcJaEtJFHU
1iBuhIKxqt6UX7NyHW8T54wuc2uT9q4FA+yV2Yu9ZHQkri4WK/R71mchTwQ4/jU1
/7qW+goZTw9lCyhHwYvP1wc5dF4ZDCxaP3Cwq6MuYBTn3/b8e0iFUVu0nJEPpo7+
N/E2CknMXyyTg9VbUifMfd0ubEDQQYy5k4DshTlugdSrnCDJS248WOxyBG7zZ4BQ
vwT36DzJdu0t/MZ2NjIQvEY4/e1lXtcjx4gzSG43TEEMw2kdIHN73kDEeu2Relss
3ca8a7yndJmytZpC/t05C/xoG0//8oq4H5+lY/eDpH4HV4nNWeiWohQqQy/D1ESM
o9yNgxzSRycivKf8Z9emtNFmELxGMYPeh7Bj35rQWOvtYMOFhZtQwTaPnouelvc4
QUK/Ng4kUcJJGO+5J9FTd1hwkErH4K7E0JaYiPq2WQHvW9vMYmzmFYlR+nLYrBy7
QmJrC6pepkBc/WDBo8MnanqxLOez//vHmak0V9mu6Pd8SHjjHLjsaqZnXWcyylja
vfFgmcF7ivE3M73GU+GSUM5xHWZ3fqygYdMww7x0zEl80m4DpvMe7bBCU3XRklSV
e/XOPpzkITj1YvTl1A0qaXWh1A1RVigCacsR3pxVjATpGrX1y4BpQBr4YrUkBR+F
96QGE/fxSEx1bKDKyGhNkA/NCAtP5f4PXOTXRhPN15KzW+feI9Oa79GNiTWkcLF9
yGLmGG4iKr2uKSQ1MVHsCT0nsTbku5ENlOZAD5bVrus4e8u8fcaKeB+qeztItnfz
6qraER2P4ipbk6lclpi3gEYeHT3SCq7byFpGQSVHYCf6etwgctnWnN3+4WGYcMxa
Y7Cs/uHSZxoxF2FAZncrNVjIUJBWICQkuLiwJ6XRuhQ631SRn6j5XmD2axaGQudE
bvtCAfEMzeidonhC98USoQJQ3vQEgqGRZvFntkhumRv1fgCu1G8gADynNw0eEiyw
WwU4sMzCwgLXp+k9VU8f4Ua9xHWXcgf9os7M+rRci9yH+8mR5WCX2bx+Ex6GTMUt
2u8+ZH9CUn25KQuY6c49lE+XD5WGfslxc5OrfG6rWJBrTGlqKCcgQl8cm/y0E6sD
6Fpl73Y3TPDnV1L8W4Ig4VUz83290orkatI6i9WA41GHDUKjAW9J+HQnXG4URgHB
mEsYMHtt4mT/7on9kLq+IwoqDzJWcqTYhAvxOWS9BLIe+E/vsxt03rebj7aBwm56
aJSlLRL+jZfH7Hq+jAfjQ5ooATm+51G/5Ij4hFdsJgOKm8m0rd8P1LFwTc8BFR4F
/MyuB5sQGURHhKl8Y6Pkk97SfK9ZyXC1Lcrf4rYeDeR6DnBdcDoP1c7wbol/RUQF
lJRQVm0Q2lW/1KAYBbhIIoQSyusOReC/UNYGYA+IOFoatZfDlZ2DhqIV5TS1KuIL
ruSUMIn5VqRbjOIa4yOg47GKzE0JRld+FSxh8/fEjH6IZuNEb47EarO9Ee7qUGH1
5Iv1Jxd2TF5TRl2/2wmK+OG2bOozkDyhqruTVsMVG8Tz2aXepfNwhHO0mYgwqOB4
mxTce/IikLNQ0Iez1hOuZzGRIj75XaVa+W5WMOmi9aZisYv/+uMXa+3oXnGeed/L
5lftxdO5N5k6BJYRJTMZsVfAYSomQAqzcYjZcj9mmf+46ysQgEzrE28kqw73kXCe
WQdrA9bHs9eZv42xAN+ve042xb6L77GyrqngAOemMA8EAsgmGlf8Vr1y0hgtqIxc
nCi2IrSBVAeuZuFIsoIdObTExtipRk/04/lwnDt/h5KwEALrq1FiNC/AQw46q5Sg
cs6C8MtrbIMayh/dIOj4AUMz6coOjoKFeYNjT0sQ3OzwNrUvMqdx16tUp8jlh/Y8
88/76q224dImDYyYWrUCd3WcDwiqVN1RBwNQNH/mAVhP9i2I/a/S0rKkftXmec7a
tkvOdCfSLRiQXhNtFCJ+pdnVRkkbv88VbSIku/QSUOZP4RdIFlY3RctJncOpw2Uv
+8Vz8gy9HtHQ5tC0ocnXGsgf/OhESiroodDKBUedf8rZask2dkqWsnoE+i6DhIt4
2RpvuVPqGvcbIH/2TwZwYt9z7PX+PAzuiGc3eROaYOBc1R06PwYSIOfa0k2agajT
0WX4yjvfViW49cqPpdbflOdZH0F+WWsFGT/RDE8dURpc90FRdewms6/H8hjpOXX8
NalL8x55ZgKkfzQfjoxYZUxxT3bkbkhynfUUiCcwnSIrEYfJHJUSEg4BV6bahplD
P0CHsG8qdXQql/6xUiuPWSyMIoD5wBgZVrL/6RapNFlyHeEYyNPDobHK80c9veMM
mV2uOgP1c33XjRMKOIvA0ZDfeQguMwmcO0cQfsDvQNsoDBnFCg6nFB1Yv88J/KtS
C3oQ6DJx6G6h2anhex5GFG48DAqr9w3oFwwfgteMPwt0tZQ+7z2QfEO9GZvDrAEc
TCCjc/FNBNSn3xSYsspjOh3U6VaSy/2tlkeD5uKUGDKfSYe5FxZDS982JrUqsDSV
eulySIpWk9R2tHEGgwzeXTpw9m+5Yig1JGf3wviEL3Kwza4iPaCrlxs4koa3meZX
B9tdRRmXItNgdJlpVLlgDC4PK9hF17B72hLBKHJuP0YGw1shxAOtNC+L0y6mkmZe
es1pH/S8ZexrNK5/K5f9HixFr9bviat552AUU/dchbiH4BJcrcT+gxXiMczBR87j
5xlepa5VV5z0xQdgoQfHqXKTlm58hK//Yl9rMUaR1RUWCtO/C/nUDew9NPSXBcfL
xUXcotfb+IVXTNtbGBsVgL24KSTL0/GHCcx4NmjI2CUEJP+SEagd0MXgRRdqoMQM
1oEwqWcclA0uspLoeiZO2ngnF6CV3ZZhNmjKw7KuyQka9+fkaioZFQUUV4ev8rSA
1h5eA6WrvwXpSFa8Wo1oVKIS2Q7bnHhbiNo8jiU8sHKsr3HqEP/SdbcR9k2KEPWB
OSjedGqIyjUij6EB6ZyTLEACkySrZEG4tdIFpHL7cr85fNnR973VpL3NB/Yo3Au+
HaOqszWoUy2lUdjwSabYI0aUvEzbfUqVeluNaAsB14BZ42Eml+Hx3TzQQQ6anMc7
ZpOr4SumdbqjPZ9wOThp5m3aN/bA6Ui1aYtOVnMvQAw4mFNwAmPMOdCl2ip0lrwK
oH+gQYHDO/BGcYB8XQOvA83/Wvi31eFqsg7RdIdm5x5oOh2UVtAQ2jqJKaZ3f767
7gKuwmFJnvJ/GJ2G8worJALvNxEaV9IIQeeL7rotwBapXC3nt840BB+sbx3WKchC
ZK1y+xMupoVye3BuL2GESNHgSRZHogbRQm+EZd/fsr/l95+C7x+j5SuUDRQA2c1E
6RbTq3aakX4FuNyXfnQ9bb4l84ea8dMN42UfOJx0peyNDcQ/k24zGoDwKE83dIj4
Nq9KDuf8hWBbfjLa4L0H9ymAYaAEcrMLl2d2UILL/haTY4u25HX9Ha/xlBf9PhHS
xCtf4ScLA2J+2NcP5WQ91s2onMin1UnDOoCpKiY1WQgN3s/BDFTMjc0a2QJFNytw
f/1kpuEE9qTONkH2sO8wxAtcjhBwlbIgzeaxuxkz6VrDXsy633RLOOG5hGfT50Hp
Dxq+tLoW9ciGns06FMObYhtYiUiI4KwfEOr+jgRaJUc5qD7npa55J2nO/q7Tgg+U
5mXIWxOcgV8EgVfLEZZux8vsDgYpumUOKfc/Xd3LGiYSgrcsmLe18pD7yCEOMaCj
pqeyLbWBN1ApgOH94LDLp0uTlCd/cJX2T8GNNM/Ftzne9zHQSKwhO1D3ljvYkfx6
3PiwXBkCljaEkD47Fv5p9u1URCRdFTHQik2oRwhX5N/NOTlh+y/cSPevPBOrXYOl
ZC5/vueSquGVgiRiFEkMbXCkRW6zsA0oPKQLhCXmxhFx4qRg4REmWITXfxkG8Q0W
6bnjHP+POiv1xNcCeDGt2jbxucguihpwUFr4ZpZKPniUg+FXZZmthrEnxMA91ZSg
GHnZ8m+t3NMp3hXdLM8vex1sNIbf38CHVmcmRd9hIJlJZq11eLL8RI5bAxuoCXl0
Ax39FQzhvkoQG4ZlMxXCq9EdeMAucUXi18+wbiyYqyUdCPDPsKIaBpEkStWw6cth
xrGP4RpgfUF4/rKgpjUjfu9pk0v66Igy5sVftN+x1PaxK7qjrl0fy+es3RPq8DlW
XP25RGu0GGN3fZN6LPXy0VV4LIaGtvJFJMIBdY8OjEm9fO0sfXhKq5+OIpYl+JQ9
P8gjy7DHHfFS5veZjjuzkaJgN/VGAiekp6D9R5WJ9UALRqTwTR1qBBu7D2ALNcIv
FG5v4xzXTvw1uCv1Ztb9QoghNi1U4KNvRMzJjhA6BEB04LHcldACxRx+10GsDGt6
BRdd/wN3drYNIcqpFP6uT2RX0kzrbktroxOWXQ1qDAXd6hQ98+S14ydijCpMBVnQ
R9FEbeUBCyLU5khjqCL4NjJbftKgwJxLUNSYzM9yZih7o81a10y8hGS+QGTkBbDB
FCRggOmy8yhI55RhR9pK0m1NaH5Wa6HT6QzSB1PQlNvbI+py13/3xvXp8/wM/67B
hxe0q97hIF1wQY2AE8Fj0n93wCqA7C096ZXP5WjuFlQw3ZvzfwCS9uJ6QfJUK3Ou
JCQJWMqxqXw8Hs2s+N8nncjuhy2TSAJVAFCJcIVend1i2V5puSrWbX7kwg15PCCn
X2Qp+sajBzwNT1Z5kkfEdJXQuq0iYSkNwAT/H1jhZVrfJCW2Db5ehhciRJL/mQ5G
91UaOA5xsrRvm906Np2j4//Q7FOicoq4x3/fONDSFdeEk+EqeqXVGUxNCnN9to9s
5jTnfNNviy0vCymTYDnEDD/nwxhvgLbd8C2FSpjcYyNKELJLGs9cZsXFL493pZcl
fSmza5hoKLW541oXN4EEmif68uyQqK+4IASRiVveWjm8pDQj2f9302EL7I3phWrN
TqGT15TWxrhb16FNVYeEmdo6tsf9GEZ+4DxGZeJ9Msb5gdvvnr2Hc02evtrvg5X9
jUy8lIMpHPy5k52uJqFuEqSoI4AtWxVAnPvZif/JRwrGHVVNde0JV2nRJUd8jUP4
8bsMqEg9YEOLS8WTMU+0McPDAuldeseEoj3Gd9rKYqiG49q+F5CywEYlJPBw3FF/
ia1JItMsx4SQgn5rGY56GEeAdvhabxlX1TyVxAYf+bWEXWyVuGWPzafOhvnlaZX0
bu96fVQ/MFGLdrYHdo8U8Y9NRfIXd8K+gUPBzWKbtR4sIVAyjWziUjeOCBkEUowc
2oNiMdXX3QZq5zJsLt7BBHZhkPMa0jHGceQBcV0I5pStq8hBuFaei+td5zp5cbfr
DUPjcrqZbzRvH5S4a0D0C8a+ooMcG+Tjo73g0aWruJ20p4sLwAjjIInKcN18H42v
mB50ieW2atL/OG2mlBy1yS1/YqYLjPUuSg48pR85nTS+/mWJ84vlqX6Kjjfbzyap
xeIei+xWivrJkEsSqgkZIOGzUATtNphf4XG2YDW/XHA8mghweeHCcz7d1FQ6Ift6
DqenisCWJpVzpY1r5PdcgT96H+CCJWn4ra7pby778T2BjFg0cZyFTaIxFvroDklK
IT84J2HCUgeocqVwdZ1YYQQ+QLxtnDPwJls0LfS0furXp4SKR2Y7IK5h9uviKZQi
NQf2NoZGHQKhjPxO0kf8U3ttLgt80NEGqESxWBK8rU8nWvmWpYQXSaCYUbwlgQgR
NrwSP8DJkn6c+y6pZcTp7/v7nk8nrM6Wy7EcZfphRiY3Xj+Wd6zriW0gNkahLNaY
0BlaL0NJM35p2fi4f6btMV5xBsCz9xtDGPVfdlAMQdj0nsIgSFoeuG64SXfAQZnQ
16278Tf16Ku0MqbbRJMdy3SHVNDkRq2mjrjiVksebsGwyxksimlTQXtm1mgBPqqP
y82naO1cqV7cU/DZmCYrFeIKosh8Ss/JWhSgvOpQdeenr136OS1ry8w4ofnCZBuy
wKEBqZhPnAd2LR16hRBHjENuoUbdWkUs5Za8Qlby+vCrfhBn7fCG4ZRdu2VVyneN
9oCxQD95dbC8gWFpVk/pQfjSB76D8psGdBPe1grwK2CwxIty7RWkqQ+eNSy0wnfC
Hh4jTiKvrOtZtXCtAJxj83//G2qBIjHxjIVyk+EdMU1X44O+dRJsA90NmWUON6IZ
FfIQTM5lo+JcB8pEJo10FU2ETxnED2t5VAhEcTv1IJo2AIpf5X4cJ6eilNTId5m+
EJZTj5ZyVfaZaA2y0hOXpg1zVoAAgJG+fEP6Nb0ApD6NN6fQn2bRXe+p8nE/VnQj
wW8Xo3zYnMKBFv1GI0X4okD3yOUwp+CTr//p+hqNqgfB4NgU/oC/xphlXAoZQqRl
kUt4tOq29hz7Sk3Y+ZbT/kJVc+4gMc7cO+b4oohnN0jj3YsbIxeLNCUcM1A2fSD2
wpLvMEp6qZXfToF53vE/i+iHFAPt1zk7V2ZZa5cp9KJnmGNgyubDLAlxd5fIPMU0
Iw+LUUq2wr8svxbNWQyaraTuHnkdJMSe1h94gUNCncujgrQ6IhJPRdVMqK06J1Gp
2q/tmAdWDa3I98t4Hl1pYP0YiIRBuQFlD12KmWBd0lGv+WCB9Y/FFc57jMNlmhvw
5ci9cuU4mkKpHyg9Vq7Pa8F1H0HikLnOWdPLpVVDDZFhMuZy18Y02jHI5g/GPTA4
7PL+++e8/zb9cS+pdYjplgTlPy5A5WtfHUiGqeIzi/hSPXWXzH6fA/a1Ai8sjyE3
qrXQbs3+bhsIgTq3wzufn1L2kCMh/PfKDNfsc/slqCvsqiwsYb15M8JQf6TcQwQv
MisgzKhpRAlCJHpQfzb6htnqGEOnjIsD5fkFOuMqcvTmXJjECJV2011elAX8KzdF
qZvFojtukGw5vvn3yosYhdZIuk7IcosIbGqw/gglomsFJ3BgZyTgOQI1Sg5Cqvjp
AjCOWuhDNlfAqvhQH3cif+WYfqvUiD10bBvz3CSA8AmzKUNgUytXLpPHLjlI6dK4
h1ZaKnrGv7vU6Z6b63dCRgQiU/zcvAbreVctQllREPBYgfGibSoNGmPn0w3uRkXS
5yYFJbxtb2GxNgVHGQ+E/82aRHdFTOvZR4+5lw/DB7NzNRN27EdlOyWN8IWVCLs8
nTN0a0bYkHPfwsHhkUm8hP5BX2bE55+NR9kxwiypsNjyhCkVQml+4Ydkihdi27Zd
hsP7/BOwJm0YjHUBwKAHIGWf/BZ/ow+TGOvgO+fSgWS2oWFQ9hGiN9I/QtaGQk7P
67BRAupZMGwqkiKbB078XZCMGWkkvZgKuZsTGO6qbrJGhBC2wDx/ZmzkseYnAyai
6k6CLeY1e/klhAF7m7XNEpo7NGvDlqiDHfT5YVzMCP73JXZqrycxhtImrNXb1DcD
YXbHte84LK3QCx4sMBamyaqZQNB1fMOigDsGk3hg/W9+uCkdaZgIpEGgMbiH+OMd
4AG/4TGwRBcw1i9Vjqtyqpp9z9zr1OhL31ak6WJ3zOBrbqA6xLY5Iky6iFUlqX1I
ZvD3VwIEmGpzso3YavDSACwZHD6iGv3YwMk0dXu3ukE/Rpn8o3dd2Z5OxRF1nQXM
8H/R1QUsFPOZIxOxRUHv0ICZlnKgHjp0EaWg0jPZGTM+pa1m54nwQrIRLp34FS9s
KgEI27H63GunQmwX5AiLD9XXx7IGiWRJsBujf6Gm8yYis7i4a8DjEH1uOeS7QCpJ
F55cWC1fWoD7LLECXyiRS6Q4Fsiv+as0lHOOPgciYphiuI7oxDbWGqVRXXA5Wlde
cZRX9aOFGE0YxykSeDTHyy7yAuuh2yXxZziywjm6OkHVAmH4ov1Wl/a592Z1i8eh
Sl1AvHj3uCVPIfXXJJtWqJTDZRxqG3y320MVa2XBuLx25TgTYkb1Y2XBWBcyUVaN
Pw2hfgpkl+GNdxqUqY9ScfwcRhUHEiciVKUDdHrppxs6mq0bvpKLl7pHH6+tAIap
dNBKzIU5Vu6MQ5+ge5GT55D/8Dc8CMDWnliUsHnB94JiLljhgSKctgbCXt0VziOJ
a96UpC8ou1b9tHjakX1diB08Cbmk/0bbGvZvCM7jRSg2qF5bPvIH+F85lZYzREeb
W1i1bhljz/5qR2q9GYyCuTCgRdwhOjYH5GvNFbAuHfIfOUrIvi/KYPZUjQR6f7Zf
yt1Qi7xVNsIiV2+sA0ahbQKqiYhXyZ+mcGmla89HP8pZbDTmlilO0MTH1xVyX6pB
HmEF664rzPDttc+gSa/KNxswObHJez/pBZPqcLRvGYNI+XjZ8mrUM9Ytorg9s6T/
kD4QVTpodd4ViU/u1VmKQyY4YZ77Qpgam88zMNnjlWULwO0NWZgAIOFWcyn+Sqk/
aeGlwzG+bpamX0LYAfNP/tDrGOyiYNxGJxhthdBbIjR8w2lCsnKV/D8WhiaAkLYZ
Jz0j1YRzJ0sMuO/sO/30pT5ZL1/DKbKNguaE8HwhU93ya/wSF/y+bLN2feDXrpaG
QM/RSKjSxElRs3CM/tlGBT5GcWHw4T36Lx0Xx6KZyHnuYRgnqsJK0jaWbIoYD+lL
3u7UwbeeHejF3elBt95EXRi6YTR6mJogLAjJ9z2mq2iyaXI5mfyaA/b9GyP7C9iK
9BMjEDfSdiSSRHpx/0gD/1YXspOdi4veHRPlPCXvBABePkNKnAjo/RdL2Yjy+Vqq
xQi075drLfEuoMe9EMLBkAg/AZNm6KItPisOg4d7PrVWASAOaVH7CntDsnZPPq+V
6f6AEcOrcWwYrc5x6+qDKGUsmUSXain25Z9Y6Vk3RmfHXNI9WHQPf6JJCzKCETgi
8mhlSAF9T0C9fZAT0662WOrmmdAcdS/tmuisWEaLdGxXUasay7gRU2kbD72+UBqw
AygnT9jy4rnIBkftxSp2Ac/wS7XQyObFu7oxfVHBrhu+KnhdObDkd/3ZWDa3Z498
s6vysfDXiGbdQ0IYVCp+5xy4yJUkWa2eX8m4t7yWnemI+KgMfYTzPmU5gJppRo3F
FgNW80CGREfdAkXx/GyVOUnon7LcQTjS+uLAGmj7FWL1361+Ut9lzXhWOA7jEEJW
iBQ93X2Q5Qq3842Pc83HbBFSrZOW6QOuAO/cUtf2Ca5eumX5kDHSjfRETOoEuzI2
mPzdW69IwowfEQL25bQU/Y6ExgEDN8ff2/ZwsRSFWQDKNLlVV3pmDQlqgZ3v6Rug
e4JhTp/IDbVuBixfRgVjjJEBiCxckDK/3W9pbrR+sh683uXkJoSb2MOy+yHpzAcm
0VY0hqzcJ6EWasUTbikTponOdvrTI6pum9FkBAuJ1RlaXXM7/iiEvOvUHuHU/XWb
sGF4SL1y+ih3DhITlFovhyDULHnnquPuopNAC12bKYhapazAVIoriFGXe66TzKco
fpXcjp9A15cZ1GV3lV00BaUSRs0KSlC00erVF2euFeo8yuF/S/EfeRnKm9ZdCXe0
4ouwxnkRyO+DYSXTlwMv9e+YEJY8slMSwUM/y4wke1IhiCy9gF6g9UGBo6v8IAaY
5Ew4F1Tosa3rs2sY/OE3JoamUPzMcJsWYdjqo/z5V9GKtXEo6znLDor//+kx+Oxf
WIrLUx18Zr3z4nveFJN/oOpMEehLrm1dAhzcbBPxOU6FQN538hDZRiEj77aC5x9d
B7mNvX5j+oGLqBkPFzEXSMgwKpBuPAHwhTO/I/uvJgF4mmj3ZXHpTKK8TFjfYU2f
jp9OJplYZS1PjEnk6TdzjsZnU/aOTONKOpdRLzJaQFv9oAsljEC8DAOJsyFWsb7E
y1zHqWP65gJM7RmVc/ri+Vvx1rDVqex/kQTLm9q+CS0247OeQDk136YRSIEvD//3
gVrcynGyL4ezNMrDuERYuEWEq4KAjY0g1ZSTCfDq/tB+/R2qlw+Jwa1ia7tLlZnQ
MwJcT/+f7EfxPZjlAFN+D9qzf7bqBiy8V5Rcn0vCuTYzjXdMOb67Q2uEJBX0SlEP
UPrV3yrHsS8OUkc76AGk1c4LVRFOJ9yFJs7spY6e+2OZ/4h8Ql5TpKiRJQ/mm5kc
pmyrHED961SgQALH5mQsaVlvAE9xTCtogE4pVkaYjw1bQcjTBAVRVEgTHHeb7/aP
eiE84iVYBBZyiub3mqFaOsk+2omIYcK/sWTVY6+yF7dQy2PXdC/JIn4kB+JUFb6V
NxHyPSZt458aL+3r54o80lpQSEGAu93zWNM8ma6o7H379ERNlpMjfneaBsDUM8ul
aY5UuYttxINvg39iC6Rc/+3p28tW5g3muamubGTKiXAZ7HvsIVonYm/Wzuy+2FTy
lAfWI7iWbHZxGM0dwU5nn2uKw3h521XjB8nCDSbF85DfuQiSvVjG10fSaYssgGWL
lcogdHH3FvSmzrd1HY6JtYIydmLA8pKQ+Mi+yrO7qI7Wj5zbyxZzVHWM8FOMiA5Q
W4c9uuh3YKmSSdSs0GIG2npMtCA63TDvlhK0Bffo3Eq0MRC34jY9cncCVA0HO5mL
uZ7MHcnhjtpbIu7su3pdzI0uvsFKtzvQsQs4Gpjtq5U13Oct3yf5BmVVYc1dHr9n
nrxptSx5tqdZ7XfkYuCMXrPmNiEAXjKdACWwUjusoUpbGHQtyILrIzDsecrg5Wb9
ttr2fSCa/4/AvFFSvg8W5phvZpEBQ+QPMN9bVS25y6MFaYWhJOXmEH+T09RFu66V
UnFMWywyEmzrY8Nthvqb6yo6CVV22LD6Mpz+rWTd+8CtXn75bZtjhViV8Bn96HTI
gIPd5Rix7CoaaUf14u+1r5/9OMs66oBTwYj9wgWjLTdL8q5e2PHkXn9/DzIQGGFI
8SAA2YbIX3NHpIOybtUwQIgQfa2frO/6MY5A2755QTFS31k+nohj/F8GRVgB+gis
c5ICflftseiCVNcFZygqyTRRpxb1cZ8RTxa3wes9rFe8PjZQAIF3k7xvQUHF84OU
COcqJ1/ydtCQj4p0vwfwcHpU7hkqSlOHpu85LAtNYdu3svq4nT8xEfVP2K1wzHr0
XEmkgMe93/hjwTAixrA0Z0Tk3sYeyY5wimBHNLJxjylKnTJxn7TCZ8g8uLlcS9s/
drjyQruMUMga9bzMsmySLWqDwT1Wtvae3FUIYWbo3u2sJ5C6Pk2bkxiPwSze++eQ
4iJxII57XLZgmnLVXUvvAntX2sFulVIopfXPfdjX25ivcYE9bn4/2whvXuafbUuF
Ul5zPOi8YmOq8onRV6Axw0tE2gOYt12Mp41yu+qn8zmk92U2eA8nw+2eQCpBqzhR
j6gpERJo/aAik+hxvfY1FZEK2kp/P6o8KzrtFRFyiokkN5BB7yEJNOx3H3G4dlkh
fv12F7HJaxjDWiEEriqUL8fzgcm8Oa5ygw/jTO/RtDXNDqINF6gNtcIMMf/JrtFh
3Dh51745SHZ3aMnDCIKgdZA+8wTrrIlZ15KDz+kCu2BMmQHYKaBUnL9axj/hnhii
tJJjgODqLrtmj2UNV+kbaeIhn3zxOYYPxcnWe9O5Z2Kp7X5/j7KfOwj/jqGiL1kL
+fgqnS7xwdI56X1oYDt4lRLRexnXdKLZbLhSW+f+1m1/h9NWdjIFJkEOC1wG8uHk
1fjfDkujPoGYP8Oj2nlRys4vvpMoAfXocj7IB2dw5RDYKOHuLD30ejUrY8/2tbM1
hTegPSG1B9bpCeZ1Dbp+OJSG165UXtorUfn7IqLuQOJYACj1OGhhhqDPhK1FLfJ6
sjoz/+uSGmLEARb6y27kl9GyuVNB6BDBd6qi4i7HBHFksVpEtaEyitheppZtcZr5
Y93NoWo/7guxpFQCQv0BJSJS5aquw00U2BJMWr69aR9Tv4nfbVW8rH0TAE37Klrr
TLJgL+WI19yoNaB8STouSUr/2EBr6mBVyFfpoXkFtExXNg69gV11h44vbU4+xHsI
i+3ezPvT5BBI8kfDGtP2bxIu0Xl3aBDk+4TFx89ZFfMhF5Hbwo5RliN9VeZNmrsf
MS6qYN+cedcqnOnqxcpv3jHfTjGzKq6+daS22CTxv3xtT+CDfP1HyQVy33VetBpz
F9thJqWKEVYdOVvf6UBu6IaguRgXFFqIzQe16/L/pqphXtlC7c0HPoAaXnEXwC2h
Y9pR1P0SO9F3iITkt1iGl81EW3AI+3s4eEdB8YZoNfCPsGISLoxPB/bwkxJQ/ixy
xBWA4vgx4UuXPMCwZe6xMrI2E4Bs0+Y9liqt9+JTjLW4lkF4meAotbVypfysbx5l
+rScMS/C3Cj7kjcX8j8mGZknwrY+KGb2mY//otoo3tZbdlEBfBsgJ1Mnu8JEkg6u
DbdQta76A7zgaQscB2kleAOfaZJ2W9wdQ8T6Vni/9poi3DB/6J+h6aUquIxQdNwr
lnjgZJWdsgKMi5kiwKfQj6zqouIKkwWS+G9CPqo/n1F3fSew6OHCR6bMNwpeCcy6
23uWcNp7ClxQqnZjSz6TVHvYS8bo3qkwUuiuwbANxyeqhAQgTdU/L0i6QXlXj+bb
rP7bARTfq86jI9k/dVdugXDiZu5VYhAd+jBvNs43Wqu30OhQRV05E/N+q7S/enuL
0hWkCKhn3OJPHxYjbNzdapWAk19ZR/NaX+uQmBHFFpFfVp2Jph/89paT3SiiVj4N
J4yltmEIMkUJtUiBf48kg11u2ZbDxJoH4zfjw4MOPtIZqrQTakp09s4suSbmLUYG
UKAAqcttAkRlD7tk9mwh33ZXs5xUbfLxvr7yJPdkwIlKo9wLCVWLQ+HMsvfUOpUM
QwL9efuLQZKpY0G39y4+Ce8YlO/sVWF0Za9HbVCOiix60ZpIxtsMIHMaMZcXnFkm
n6Q+A9q/m+QzMAfGX9EL88WRyvscDTHFNZt8WFKoISZhlw7zvbSq9vL2Kolk+PJp
Xb6dWp40PsbpYyW++fGHVeJkt3J4Y5SXJCf1iDJx9Pe1QIMYVBAFDSP4heKnva+l
u1uuKG5/OpZLP3ivDHD32lOFuK/NUcJpmYZxcvL9A4yhlMyapBoNkalBM+V+CFOw
CvY/tccGwPEo3tFp3/IzMyxp8/ONYAiOOlKc7hKwTvQfwZ2fo/O3L2+rtV/WgZnw
vYv0KxM1aQqSBENfFtELCaXrBfsNcwy8t5vIZzsyq6PAVwj8zfXk0vkBaNZXd8X+
07hKzwa6OkJARBM9iM4onw68VZbfCptyw+7E0fecBIzznp/U/r4YfgKHo7TA2EVX
eoMTom/9DYEUTjIy7aMzklI0bdmwM7UrPxthvSXGLWt3JR4QDKeAX/4f9oI9kmwP
9oL1zY+5KQAH/GLmKSX/qgG4HClhv5ECtQqAghIUkF13CiwcpBcoB+TJV2Q/GYmS
JiCa1zMuOC07AaHOYA882ix36N6IH9r+dQhUvLXe1AUgoOCV83+hmdDJiFgClxyk
GB1wfDc3oeK/a2TyDLV/Ty272tyQSn65d0F9tAdglpowp687Qb4HLIi7mG/c0NwY
Wqh1EzM4qZqvEHPjoUyRJWNsF0ArrNWeVDok7h+rsQP5Y22jbKlteik/MmNfwTTl
kIazK+mhawp5sqLmqeAN4Il7BXxfUI8o4Omm0aFEzJAOyafzO22Yf32nXYFoTspu
qnPCWYxxSK4sgwrijXw8E0CfNUvEkzVSYPxhBb7/iYNfDHvIRkQpOGQa1Ahlzq+e
Xt3mXAv/JLIJkKcOgh+Z8hfQjl7t99e9ByB/6ynsky3xAkw1N0mc3442ndoxv016
gYgvLKROvjls5tT2pvcHZ5xi350QTF9QnHgyhuYvVxQf+UEKk13FuCgyio3DPrsd
pHuk03lKJsE8vOEW7cd9pmw7yVDsKrusfK5yT5APLdc5B9e8NQV4nhxBBGpv2q1d
J2/tS6w/fStPdL0CvUZmLFTwDqCgBSyqgInbjRvimDcLI8QD3n2ib2oVoBctt8y5
OWfMvAMBYPlJxcmBFwgQfIajPP9wocT9KdCYFyeyj4YPv4wfXIXzDBLzbsJBVqdw
Ar8sAvw26TleXgNSUCF2sto6pvly5AxYAbiszT9jq66SguOdla+dpoRpy5cY3PXM
tsbqL8fhBaHGKGcuANSdpcm337AoPaPiM2mocwFYBtTSPlLW2GlPTVim+TDWgPkn
N2qwFi41MOS+CRFTQJ82xNKruBU8eu3xTJKL9iRP6DlzrqJpTENaOmR2y5DCoJIv
76lGf8hgUdgFCAI1QfCgBr9bV9c7TKnO+8lQJTN97CEWoOwq+KbpKjFB2TaM5xoR
jy4wrP0HagQ9eN1qYlc6qprUCAdwKcnE3VmKztsp2uubNYdLLiCJJcLBII1Drhu6
N5PClra/XOqbz2aEAhi+J5c6cNZXAMEMriXThKpsS1WKyWf7aMJdGocWq08e0kqw
bdnXY2qKbUj69CBxDVXSt5gh3uhT2MR3M2kxjAomzaxwgv7qVHC96pnnJEYeOCda
YwHrgK0LlwkMEOzDcTna6uW5ZOZN2LsSD98aR/4f16TEJVv3U65oZH4L/Ik5h4Le
AC0izqhFfsLuiiGDLrXLPx6GhTPMbTctE9skwuinBpyiWJ83yiVq9giCBR+aS75/
vMJOyJTjIptyXw5S+o627J/yE9JJRT/8928box3AdGU7Db66irkm5PIl/4RKiP4c
Lt20XbLTiKI0VfyCEe/A/W+9NLBEPdqpWA5DpG35MaLDAiRbKwZOAZ5eko4lHPt9
CGsu6gT9Ewci54VbA4XR6a6bEeqiLRDD5DNQcwMwhPx4o7tF2m/OdVx2+VnWTa9p
w1fbm6MtoJzDRhzmOord2QlH+TXVM1e67lIUwWTqZqgmB0PIxKKMd40FsoIjKadI
JQSdNc+O3bWNmRvXtWfBeCiDJDio347dFl9eWkbxSf65jFFLmzVn4dOHtm4gViVd
B7fUjsn562ZNIMWqqj14tUJekSuAIWghelk1/dWZBvFJFFRKy8EVVz01Oeyy00pr
JM1d2lNE0D5eY0C5BPWQKrpWMolgvjnDfSs4cMYoM0ZIyanBeYJJBNgprMI1fak8
sMKgYg8WlrbcN6cJw1n61pWWuApkecieQ3+AbTX9TLA1OASlzMnzj4+WR8yzT+S2
fB9Qv0gHPfqXrtlfrBJBHaA1lNDGwv1APYAQ/c+UMqXgdwz9QQyc8KMJnZqLD4Au
Y8xhHTos39VVsntOJBlbQb+7YmrOZXwP8gLCorBIc6B9kA7ppRSPfn+n2tTUlwTG
NyJmdr856GztSUeMQ2Xy3UmAbbJLMy3ZLEfC6lTrdNC14bIKY8mpuB7XlzFtOGAG
UJD+9gvkWD5ROmAxNzIoK3qVn1vkvZCj82GYUteXQEB5hcX4DmwBhTsTXt193PaG
w+iSptWMl4u6T/sOoQd0ocoTprEhyHK0YoNJqXXH2ZmbsxJOksnqVdEValwp7Whh
8xjz1Kcg8i42xsZHwg5H+Aj0uWd102P/frR0gL2kVyHyO+gT4Gdg81d2OfVHdqZZ
GhmadH18TfjObW8e3u5M27YuwuTD3RKilZMCJEQeiX+ZvqG3uv52d3DOofQoL/Qx
Duhwhx5NMEVrwiMnocTXJLsyM2yxuF8UJHNl7u1ev25l68t/3o94KEE54wGO+7Yb
1Uwrdi+YfxkLaDAIpGWh0xF63vtHLaUYKzGxHOd+kAy7aFLfTqpl4YbdrY5jcqCf
E1NSOgMqvbl+bXIyU6XXm6dFjjzA12xtEBMGWM+EE/g67Z5yUmQIJUslIuF6evGn
i6dhJ63VdDK6Ab/m6zfBmhMKWKDjCYTKLhlcU/Fm8DtPVBUyRGB6/yJ02NpGuu+5
dLO9oU75hK7J9D5/xjhgCc6CklLFtj5ZXbiIHe7aLCDvwHJeLJoHvCbKYSYzp1HJ
aN4+G1bzGdFTp65J7ZrsRRF8YRW+f377bviR/yuRi/TkrnFT9ZslvxgDi2DOEblc
BGbgiHoJ5xyaBFAZDYUGyMYAMoSUJgB//tck48XaXqSpNzFGfayuuWWbZm+EV6yw
XUCWqC3ze4dQ68+pX92z204twRT765llT8E5UnL3ONLU5qumzOnnITNpQguey0cT
4jlM8QILoJ1hiztZbPjyVFnRKVFjiccdRz2U/OL2lbe/S8CtBNRV4t1fPzFGMnZx
WmrcA9kDE6Wh6B4a0vO8rE36BqixBz2NYVxV9o7EM1IGDuR3Xl9lLGfIL/JSXM1a
yxSq/vcDkpgxN559y0MIm3Vy+swIZWhk2ztD43B6e2BD78Epw9CJSdT1gsQ30j/V
IYr5sB4JUjHKRrdUeTDo5W5IuZzeMqQFY9rkDWYREii2j1wfUX6Df+n0LxGvZvTV
jwKYPIIHXOkW9xYfEaT0RbbYzjsuvthljQEd+XrEeyk1fdWdQNI7OPeYii2HFcV5
RZMkp1RnGJLQ0gt3mFKt+4WI5Ilg+erFW4eTehiV+cyACfLifVhLr4GQjGQpyymP
jRwnXrhaMTZFR47sqq3QswYzghHasHfl5au94ZOjBr/ahvGTDJ6vGA9lnZeIp2FP
I3ljXkL6eAZedj7L2YoHnbhUn2h6Lmd7wAwLx8ut4dQErwFSq6T8juRPLOhdT1fT
HBefTs8TtrnR7vQbwZZ0FuHPOEGbd+o/XPwZQpE9pyALop6IJbDRE7QPaXiVMEd1
c9bdvjSKnWXf4u6Rc0Pg5+tO2ELTTHuIcRWBa+koRjTNDjpWtoU4+076Tw4va3EN
vFZsjyBJCzbKFhLf+qpaPXz1qH3MyW11uvCI4qEOc9C5kS1p3nl82o8wpHEL5Aw4
xZK333jYbCWfVN5JHNy9RzNEA9efLAU0DDlQGKdVXxDDMNVAP3oAKvqHJtmOK+RM
ZNFr9ozpQs+DMAaHYK3TeJ88/1vrTngUMkpUiDeQvl5nENQYB+BxRGCgNTr7+1CO
EXsOj2AZt9eYxFiCRHqfbi5v+FxtZ41AFW0LtyPattHo4259cBT8LNEMYogXtiBn
YoSp1TbwQRxc3hg/jt82PAB6gHQNKkFmaaqs4O3V81vYhhiQbuhEYFUgjq8b0OVX
5KNoxc6Pfe4trqQ51XEQwXLgw+4xQJ5KH3n8h0VZKuJ0P1Dw9J1d0IUz4KP56ylz
hNIS/5xj4jePLLzXzOD/UtRhCOdgO++uT8FlNhsLVVHAUtCYjGfbDVJ85DIO6Qts
UET8GMo4t9SBvn+P3T2kUiU67LJL2zMP6qda3hFK4V0b3nK3qvEHJNXdTmPKpvXO
6sY/AwEmK/HxRQAAz8C6C9mzKGEjWGcSsbb4iTHs5RdHKoR0LBi7defYXr3iAwDN
dMukRgc83GG+PluYXcpdL7fNdZpUkPppHSiLpP3mXg902gHBI311NMWYlZiSc0Bq
ouZUOPzJyOtxQo3HlzYUlURmHQbFrb5hbtBpPsfBzQfMzfGUXeXG25qWjSOUN9BU
Kd+3Fj4KTcDtUPg9r83AOG4yMLl9NNPUhJL304t6KwhF6+pnkV9x7jN73ruoAZ14
UmneFMhCsVjEZWROmI6dleQtSohp/8z4/ZywGPVTFrfJ6FJMLCIOUvyiJUjR7KmA
d1cncGRET6OEKWz/dLmyakybpJOfGQZBDMmSKM6oGLYo2GJygIZPm9zemLBG7OS0
UE0UiLOWFOzZbRL9XAlHm97elVTIpoMnmYC3wZHTRbvw1mqPkgSTM/Tu9XXOgbwL
R1orhW9iddzFXAoXQcAkyjXNsfWvUNiXTtkbfapt3uEc8HEWqTgK9t2WueNhQaMQ
mBTyT2jWkuRRvyIp3v+rSd8H4MUPcTDwcqZmjGOJnI8OP6VIcj2tE3WyaAgW9dFr
/VNwcdtzE/9WF8OxTv0YC6E+uNk572Fc9hbbbtmeDQ4xBBLnefhy2J46YbHgliNj
h/LDsWfz42IE0kdXNDcBtXtmr1JbRpFdzl7gWOkzRhtfzQ53GwvxwKEtuGorqzyk
upMNYC3VujBWa9nrruAuJHkbdk1Rr9Jvw1qv4c+nMEM=
`protect end_protected
