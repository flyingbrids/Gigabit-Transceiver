`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Ihok7v1T8NKnYDVBwq+Vfjsmk2T718vKSBJ+o7hn52cbxK9blw5Gd5IkIg7SljZU
0knSkQSm5SrIfQE08/ThNcQqIgkw2YgsZhBkDAYrO3VQbE/l4Y0/CGrq8CzNvZqS
l1kPSHerBTFRq81mePex5XbYVDlQ+s2hgFi+DGyd81SnEvHN9S2TW7yiLnaYSP6c
lwJHP3yvhs5B0VK+F+7ye8/uClBk6qOKUKUET9ND+eZukZO/7rhizwx4lMn2SfGL
HybGbC623eqLMX8Q+ZfYL+1y5gjHBJnI5TKHCvv0U4XgJcnaSBBm2MfskXq5F8HV
7413ystWGgzl+yCs07OLTA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
tTADl70QBbyyfGOdIVOd2zl9AGOfcTSgeFO+sPqFjeXW2zoZZe1ioWDrjQCORrTB
6xVOVZ4RVbJXSktToD95JbvZFEbsteKmi0gFTx36aWzPKXMlrjaYoZVHg4n6EXmC
0mhu5PodPIK8oTL/hTT3b6T6PEaytbA+/QxiGsZ7JNk=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17488 )
`protect data_block
gLKZUNXLak614ex3twxTGOQLTEaI1m9tulolQO+53pXFtLjNnJHzIupddOjIGSDh
5PRHRLf9pfqKdMceeCCG+I2yGji1UaqKwkXE7D6uFi84CvXtp5SutDVeq9tUhDGv
KUMHI7PD13CDdpZYfRY3tsNUObdoJTdurb1kIftEQSQecltThn5Ic/GdQwWmUYoi
ifTTFn0N6AzwAGXpatgZwlArIWCAh4fwm2fEx3mMD1OgkMm2j9N0c4qw81Vw4mCu
aWxCF9A8ks0AljLEUTrMtFuSIcLPPVli8iU0JKMei9x+KPu6BnJo9UPqHwxjF8R3
DtrCbaIcTp9D7KnYCI4D+SPk9c4v4vkCNTdFJLqhthoThnN+Pj8DKWwAmou8vDQr
SDmTbTP6nti8NgscdCRIRXbqz4IwKrUES16cGhcJ+A8hKvGkTEbOew8i4c8VQKkY
JX/0fEJk4ENC1J1lmCyw+N0SpHoHT0RxsbOTjLW6TWxsenwBYcEXkTOT0iG15bf7
X2BgGFJ1cAlLEdo8bRFvj+JscCLHfRygGTKOQTZ3Q+Cgg0so4NBfuyv7ok2pz7mP
5VZeoYqiS02iiuoVtV5gYnawxBo4/Eb+uhoUIJASa4IjhjtE69fAvucDpKr1kS8W
9Z7w9nQWPJlTw/vQ2zhnoganPoMRZtUQXNUcdOEyOO3fGUEWyzive+jbJ6pRT3nf
EUy+EODcBzvQEmelHAZJ2EWCq53SBxsIvgWOQfUn51E6qyz2BEZ9YgLD7AfmBD63
yg0cmFciVEVftwqfY2r3E72pwaVPOe2qD9FVj+3fSq0j089+lOZ5cMmamnF9pGwz
BGt8AyVgrrltGT9mQ4ColX6451Czxar9eRL6ug4dnirgF1jFm3C+xMamzarH0Si8
s8YV7HaexS3dSGrM5vk9amiPdrtZ2Kzs+rTHQmBY3RoNrPVWeKibU9JcEau9yziX
M6oQn8KZffEic/OgS+vwfliArD/mo7PRbNKsZisMsejjV0Rj0BoB08JYBPvCpQgz
KazCVV+t3Hnx9bMIgVY836aPRTicvwPQUF9JmWj14/FB9WnpdTRiGDvW+ZxXJfa+
RIPbTWsrG+02hKM4oqMFI+05hVGq0mbEDWE2iygX2TSmEaF8IZZGbPALxIgk7hqM
85qUbQIqfONY3OWWOjN9WSX6B6XoT161Ugb2iC9SNFIV3Dl/ydjdIBhVYO6yDKn7
T2BdJ2fBo9W/sEKHe0S4NtiGLh9b0X6ojTlROV3M3DJN3PUMx9UyIkhhOXfJGDFH
y5bB57HHQgc1Y0yEuMODM2Iw1twJ+9yHtXcnJYYXe6yWHZdNK42GIxPdTMspjFgS
JuvlnB6leNPNYqwRxAz0ErnEWFtpgsgaRv5rXYLTq0RPAttJq0OsKkrqbELrJp/3
yL/qV4kqRPoJW4dVqxHEb8RMujMavRF0zXUYN9JYKzYlBuXkkbfWbZQbv5xty/02
/1cCiliXTXuvroMkeXPlWBvmiYUELLTZ6b/DfP7GBW+KkRni65XLB5T9ntsAAEq6
Csxmyn2KXX4tlPRScNyl5Ynx6/MfB7UCxBs0pCfob99BJ+DZNr1MG78nFT159ddT
AZlIaTOpZFdshTV+oUeEovJM5amC2KMUDI2lSXesuJ5Dl6m1n+MSSLE0hcMDRFWV
T1I++KTl0VYVJtlvIIXi0wR90yA2mglIynIJZeVNFKUrnqqhiQMw/6IbGx9H5+oZ
oakeBzgUNa35BxFdYqvaGAOu+QIeOYPy837EfvCUhTzGYuKnjDxaNprJa7BTmhBU
qsPEAF1Jged1qsLhjBTFOkvP+VPCRyufdVBj10kb8SViLb7lbXL4MOkO8KqbAtf8
XMqRvInSc088orjnc0/mOOwDUQWBPKeqX2ZbtRim4QUqsiQz/RY4XpqksvLoRLUw
N0TihMrj94TWcKOk0KmlD1U488Rn4kMtg050QIjmeeY7u0c3c1AeAhr4zQvgoaIs
5SVz4bCH9QjuyPGNbMWjO6CygxL63+2hTH5ngzepVpFg4l2TjRro3g3Lm46OXraK
xH7r8omeVmSwMaFcjyKXUQlTo3Labpi4ZaiuzXqchbB5x6jnbMvJ7VP2Q1LzZdrj
JWG8Gj1SGXAMoZPRJ6TMJ9P5As249DrQ3p/ZiLXz9d1KhOB9QrxppoMAJfWc5G6g
wfRdVNhq+Cf4z1ZNgFrw/3a2OGXqVmJI7vkVKjl9adncnYFblQauNubHNPhJBG8T
Yuxk1um2YIhq48Pl2JoJ1RO3KIi7b2luIxbU1ax+5UhrQoEwLXm+Jg0hHihF9aoi
6LyEE5Xqg7j+N0Z3YW4VXWrGqdo4AgKC8FVeYRaLCjQ1F8/cZpXmJXZaj5sUJTr9
WcubsHyMG6BYaJIlpk4JlR95yKthqbXI4GOkp4LXiWvC6PDHtC1C5McNcu1byvQX
uZWedIk/D4n2xXv3iOqZEMS4wdhy0TNn/5I9Z237pdzAzk8nr8IZCNYZYAiI4Yxq
/WOm9irCj8GkihBya/aILfxCPJlnR514v0chyYSy+qExdVexoGwrOUPli3du2fDB
0AFkFD4puOxgGOyJyElFDAOMfLwa0p47E3lMalkLR72orITpJCzT19lYeD+sNKO/
vWLGsmWIzL+v79BxHYqL2XQUp856V0ghDqiIBplg+jh/uTUNhhuzZBnt7BaD6vfV
IG1Uof5pSDjvfj9SUGZT9D9viKikViAU/Nsgud2RmlL8MWfcgrXzUtNnXAzgx/ua
8KKJ5IkPk4UELl4wOTbo5hAJLFCaNW+eD3D6Ao7YX4uTQI6VXAjyQk8S7LXHAcfR
7d7ZdC32KRmBphV568uhPMRiq1UrL/EJCcrAe3+/ycXiycF1O0b+QE6QsfEtv69y
HBjKzegLcZpIniHVvD98qYC+FjBSEcMYwKSZqe2WpWm4JnWLNWh2wwUOSv2ng/cf
diU7z5xotwoRs3XEFWhbcrBROorn9rXt8IzgnJt8zZTXoHUAdCkxm2DUQHwip5XF
o3OitpLRSl1JDUwoe74n3igej/QbQ6xABwCI/PoA5+hBE2ic4I9QOOklAERiKhWC
nBUUlfywbIF4cEsxT9tWRlghJhpHevOzUM9NILhGD/0wTmnM3F/cEdgwKwbeIB8j
2KDBJWHua9WZ/qsUo/1xuA1HaaibokC2FXMUYPwf//PtgxSOoeU37ibBXq7JNkqh
lSZts7blqsxdc7ENszO8kEmjDWraTkOXNCfmKAfmX5MyQbVq+UdFm2Qgc6tHvpb1
bLFlqQEwBP4CNbbzO4lnBIOvNoXr+T85DoJmlO08638JPsaFskst6rCvBU/CyKSS
XwbS5CG5OGNI04uF1xhOI4CWxo9f51iUqAss50nVJ3ix723eWBY1nivtYUZSoJFh
PFfRxA+HWm5Jea7JzvlLn8vGIEJ4IMeD9+Ou7YFLX1k2DyhNjw4kj+cSxgo7Qchs
PHS3O3pVfuLII4AdNKCaZj4p0F8VjaQ39yqWSq+oQiJuSEOMneki+LVDvo/EQ3ny
NZSimnLPnwyibWk8nHlf56YNm7SEicqbXy7P6r9+fsEAdIQtL8V0A8sCyiyE80Hz
FJDpd2YoxW2Bd0KNJ8gnzVcikzh+e2yHcHwbIt720dMvF9XppGTvJwm68Yv4k+Tu
xK7Zz95DyVqvQUFvHvA3VfGwroyXo6StrHEwNUFaspPShW0c/h2I4ILPjqQziUm/
OOvYwkYFhoZEyceOC34tV+bgaou0n+A61zQUtitPL1AzVi8CzjjG9+SAco28ke7g
xtjArOg2mfcz5iaWk4IXe2pqNjW49TXi1IRj5o64tNw1+EadGIrir2LU7bwR3nyg
Vzq3xY8KHADIZnAmmjACE6czNSP48FZvyJQ2wJxi41O91c7yO2Wywtg9TPYGMyAL
Zaz2I7ZO60OA2eLDLutAqgUt1IMH993XZDybW/02dOLxFzxL3nqm0uw1SD7m5red
CMKaIb+7SuAehdggtCoW91WqBQ5i14N0ODOg02ceSn2rDgdYQVpbCBV3/vaI9vxM
TZaIwPZQWgffTl7cpe44RMEMQClP4nzYM/AtgV0QjdJXfqh8gx+n2Zmou+OL7JmX
S8wU7f7tfbUxvdGPLDsCtNAja6/nwt+F+ITkX3K3GbEF7CSxWggqrUOQ0HxWWMzh
OfanlQXLZ/AnczLNmdSO51RmiNEAx0W/bqYKLGynKBoGZ4OLOTPoEYlMwFXZlbZo
Du8+33C7IhV25Ew9pfsMcU/rCrYr6Y+xCYtSa6gHYJuAF6hBfR2pFjKCcs0c0N1r
YuJFpREEXuzx2haSvIpFVqYtRYBySu64EUB6VqxRaiKrOiBDAg51JMfvg2cLUwku
r+F40/fOFHs605MLBsZGw32YlWVtM4fJqRdm2q8fRbGgXHO/GXpqBX54jdZAueOk
4vTnqQEbhlHLb0PXekoXgnziuZrzt1UjkmQ6KUDyFprDB2kO2fFEpQAWERb2TUPm
K6rFMRfyNM+kxm4GbVmQ6PJpjBYukGXRymMp5GsnzIaS/guVDWvHzYSChUTnsTor
Dw0WRWHHItqH+XHx4uH2B21dEpOr6APYNYCQfG7E/+yTB5AZHCE0e6J4+vKVPjmj
2hfsRA+MgZNtLmGAVxZRjpnAJW/WKaQF0PRZ83DiNv3HeRZ34Z7Wjs8wbIrebhj2
ho94/9WI884439L9SuoSv7AOcgqUZ5mbHL1xdBV/bQ9E843fc/s0xHDvd1JD6NYs
auFznE+2Wg9q2fo7cNyHtxtlvoq435nod501DY8h5DFa9oAFnSVcXU1VR3xq8/Ft
4C4hHyNbbh+WBZT0z0zyS5/3d5DTpFIKTPpokyl7SW+J7acaHut8pRx1MH4QQRIU
liUkXkI8voMWjt/lNxU2e80P1MaN/vYEsthpTPT0LldYFlGsNeHlbzOLbFIdKXvm
DkQr49K22jn2E2SqQIq9Gm3RgVh2iqo+nzbupY5UGbtxp3v3NotYRWT8myOnvBh1
y8IUCnK7EXduO1SYer8bKXtoVLM96eAyMUhYvOHTVtlue3mTb3zzC8fGg/K9mQp5
+ONc9RJKILucXDDNHmg58FknxQGWSbyk+O3ckO4uNUXwZNYPjo7MlCiyYGo+y2jw
2VFPNQlRHMmZppnlVuZuQz++pK+DmuRSu61HX9dOcqSknJsjJ3c6dMUUc6f71CuY
GeCVh5iKv6eSopN9I2hPCmcjF3VQUkELp9v2xMQz0kehUD7Z7fPNe7jF1G/I0/+m
SW9acQvSOmoeb+99BK6EetqcmzJCqrEl2LyQkjylq6OztE/nQHcQfJmjnnN38htA
x9df9LAlXypfqgM8mHGNpQcPn/BNdExfudX2URnUjDfGnlUR0/NCS03ueKjWGzPP
/iapTdGbu85jouaHCGMnwYGq/h2hQ8IBocw6E6x0chbJy1VJgOr53eebgblXkLTF
ibIdpIHhLleQBRxsrKXFWPprlL2yUMNAqafEXDMZ9VDzgkw6M1JEPUlwVi/9JgLR
0+Bw/t/NlPGNztOs+Kb7YgvAyauOshKjYw9hMQ+lr+jPJgw4eFZrLfXLK+e7zJ+6
tPYETAG0hC9npdC+m2h4wp0GQErtRCDnwTvRk+5AjpQfJT/gEjFACIsVPF8HPRML
vCGVM/qFlyTqdugf1h0WKN5nDTPKzXjKhVhKf73NrVPOI05X7rjex9y63vVkBNqv
maKx+3wgYgAaQJR8PADNdMdRhlqq+/ZpTORq5HcX0vmyQkFk99BKc5B1IPJjM8Xm
GMoOgU8Sxwt2aAR4GpvTwuY/slF7bhYT5BdIIWOoOgXVXrmwdlYafpGJPPJAz4nZ
wXo4tChMGfGuID72fbqqlADy4dd4wgd6wuPd9+l+WLs5TXQqlqRHT/TnRNSDVLwY
B2RiCQsV7TXPOCOe0dhC9+XPDkvz288RgZ8nCTyUntDoJNfBHef+0hyV9Jmh2l3i
S1fmJrRIoPTPU51RFAXgIe6qVDjn7ieAssFmWlbHWkZuo9MvOYA1Lii2TCmDQiJd
5ExCbYKuupUvlAGApPVJHvNedRE9zrTKRlLskNvgSrWZlxsKFfKPscyiuX6m7tHv
IKF4csrhGyJwhY7oP1Qrw0UMYABpSqqBMzHbBYHPa7uSLIDHW/6rkwNMt7N3faEp
nFkGQSK6i+wmgQUdhd34uVVk19GRvjZCFePVsxBhwv4b2NlErCl3DfAHJY9hXK0L
G9et8jpfEEZsqJ33uYtAEnJabW4kZP29Y0dcbDSeTwzc/H3tszkCVk5QGjwK3c7b
hfM/afw38Sl2wzBrjzoUzqj5suIlcW7qeBfZ321MrfBtukfH7092k3WW4W3KDvtL
immFIgyhaf0zO1Im2VtOpuzTu61jAUQlYEGLwuc3Wk+07ivpUoSEHddvTMG+gwq9
BzNQaKfzAo3B8GPmbDecm9c47Q7WgIyYXSHTPc1DSXoOJnGK4543J3EN9DKGetsQ
s7UakTaSqp3hORtr9K8/3pYIvwaXHtffaaiGEV5Y10WPHdiQxyCqxIBNrfZEg5wz
ntAKDDQthlASOqDIZ02Y5GbyYIvYY/TNG0uCwvnSmtz0G4iaa23pwe0IxRViCadn
w7OIO9NRa5eXvzpAuSHrMhxCgh5DaCesLqffC5ps6YMaHfFhvl4vZVOEpAcD3uZV
BveiWuQS4S9XSBoo07Hu0Gdvk2e05xR/APIJ7RS1bi1H3W9/4L/vFPUKqEEyC4kS
EkuigeRZ8gAdNvsIvSXPyQ3c2ZwCzVvq+WwhCzUnYEdQcimRH9A9cjIFyHgA7CMK
n4UMCkk/0Xut4NnA9TIjWq0X+uEyITF7xwpYfwbG1NlEP/yJdCMtgLbtpXF65IM/
o9ysLu95MXw+TIW2OG61SXRPQhuq/w1GWxIHVPAbz3MJ5wptqfIjQS9KxU3RtpGb
IzgZI922p8oVjZEjjgNHyq1zLpeprWwl+WB2dz5QpBWgT7N8+0KtpUcEkaH0MUDl
MgpLDKYqLTOg4x27JTpbymXHD7zKdEeX+cfLHBM2dGzgmHnsR/o2Z9OA3rVc5AuV
3vNCz5NBO3HlL86y/8wAP41Lpmcb9eQZced7iiw75nmxS/cJuggTnf1gMpBFKheK
9O/2CuNYd+eNG15QT0xal28XCuOAw/EAofO6WpgR26EwyHXMFn/+yMlY6phVrcc0
YT0ZY0dChfDbQv/+wPOLRqnOlJgaQnMm7dYnMqrZN7khICj/UzDtEMAvyD5KIbvr
JcXog76WyWhEz/ZCgfQ7IK6k2cCCqWZ4E392vckIoZVfbzzvK2qBP5gK+vJuUdav
LUMtjmVXHptTdKPdNyTHigmJF65q034NgK+WpXm7OjcsfpvZi2jLXPm0yzQo4Yiw
xnB/OPL82p2rUgcEq6Gt0JuBJs5szzInIF13PdoD/6wznbhA6eFVNlb6ieIKq1Kk
b4gJvKtfiO/1UFCL37G/QL6s2tUZ4uUCzqwre6Fiwk7lEdi+9nKngOVZrie1L+Sr
9U9hd4SVDR0jAccga2MxrHh0MNxPWwYBXqtfqa28NTSNq/om+BRHZLk7IwUW/n2q
RVUYLI5klEIKr6puTpzUK/gOXQaj7qHVFLqrOhiV5X6ZqYmOoW70T98MYDZcftZq
cxOQcbmATT9pxDgR6QkUAP/Fl99MiD8QWSO+7cFp4CWWNMAVTWtUo1D05pM7NKpM
uiEvgILYSw1YE2K2lD9UQZvDPU4Wy35ftrc3wC8544iNV7TcF1ZwvkSQM+DmT+6o
aHbYxb/fPSLeZ1xdXHJCPE7T3143nDnGIYhC/5C+HsllpPodKn3bGnry3sfXn6x3
lFot+Xos5HGFIoY0DUxCfpicDJEXcfsFCiqkPJDjVYe4p55WL8Dd7TWcljH+euMq
TOq7HdTo2xxvMXS/yVpgJbUIf6/NR3VNzSBWcEhVHA7sLNFLUaYgsgGd3YisM7fS
Uk40T1cW1tNPVDhlqcbyi3Qojt74++5CZASjN6zEG20k6H4xk6Ry83QW5h2+45ZK
e/b6+R7eMnTVH4bEGO9YhqqUZib2oUkz0M95c06s/O4pAauYPJqUiygzV4R9gkx2
OTUT0ueCKYDt/pSeTPO9hA1XfnsKVEKwVD+LQbnKbb+19u3zBNyG2xf4hSkVWygc
QOSRcClLzHou5FXi/VFFrcX3mmRSNo/3NlsCsstm4W5n6IQd8VRGMBaKuqQUlZGV
OJOAxmD+C5AIL5cQQEuW+iK9FLJculvljVSQzQzT7p6D1d3FcwwbNUL3weFJFJTI
RQzVhdpHW7Fs9G01VjXQiMr5/1TcX4dmaMmw5hMDi5m0aWqzcKCuH9NGHa9UD01c
/Q5CrYVoMoaR48rQLEZZqzEtsfbEQQ6EmxNSGhsU+I/gjm+dlviYVA3oWNBevaHX
b/1obkFq53djDgDCQid+g/KWHo/lfXFuinQH1fpaR8e3sDd6UIBsU/vMmTgFDGVO
ouTNGQk67mZrJr0O0xyD8fE7WaFO5BUVU46xHKj/3VkaDP19fUkpWWF3267Nh0q0
/bhgTHUkHL4mUPo50hhF6ka1JcKHiDtooiNfYUxdxkociA1XcCQyxZOrazfpn+e0
ZaNte8qtSXLl1+RZpAMLr9axbFviyil/a+EmK4GKSdXM+EtbTNWdgZ5xBCfvkLr6
R/kEjwm+Lk07kqsBBEGYr4PZQ1uISYIaSxqzbZZMtnYDvv9BL1U0n4CNkiJi9MOn
SFLUkbwnpsHWHMQVMHI/jrlotpfH1feb0/yOWNGMI7GH+3SrC9CtbuQA5kP+2usD
cnuQMSmIiuOkhafnQosODvuGAvFrBI+GrOjnrS8oqRmuI5cfix7ejMazISpzDG5O
trxE4yC1JK3RARfSYiTQZ2HvkXdQSuHaWBhdc4sW5m/hfs9ciwnshuYiWOz1gEuQ
lQtO9GCQWyJf+nqC/WQTdAppRQKkww001ouDufoDMaG35q31TF1byyKQR8Hg8poq
jaZxKU0SEaeHCCn3DO+j6Ay+6OURNTeDQeZDDQBUsVI/yforfrHxPafIhU6poNAm
6RVVbhdwU2Mo/dfcHs/1P4IxpfmZPB2iG0kYYHFtOdTm4dOwSYjfpMkaYVekojv+
5Tf6U4RQY6600Qi0f0qovU7W4h0R0D+qtJFIz3jZqshMcvOS7ESEyDdCp3aSr877
4JOnCEA2GadrwGwCpniY77HdBm25TmAQG9st8gfXJPEYuUvUwsA0kpPBE3Vm2JPi
Cjur0/VaIwWSa2qzDN5GazJKhHXbuq+M3WqoI/R6DtBccp/GgxZvd5qVk89+LgZo
P22EnS7Sp5r4lAQiX3rWFGCkUNP/X9ucrEatfwTuro6cI26Vjd3jeB0PzM6i6BuY
AdJ0Yt/ay2izUvepfXGOkGfLNYqe4QBqjIDgLyPc1pVAfr5iFt2PDAnEdegCJlvB
LTCfs0+8hnSW9rM0/Fq1ofiNu+rtCSP1XMcHD3Fuur3D0SLO/Cx9hkVbL6OWnXQ0
fo39JcvimBga7sFJ8dAv6VqN3ec/6WL0xD2UKifw9BJPUAZ/8Wp6jn0DuqZ509Jl
TD8hIIQzXeX+sqQBFFe0q7Irt7PC6CSvH7dDrpDWErUDVPD+WW+ni8dnARFasTYy
CCboKiF6m4XqdNgB4tTsufwI3hu6GrNWE2Nya1c/s05MPzzPnyggpwCf66quqRM3
I3zHHLi+Twd78vJnLWwTOP6kvhEqiE258M+XIVRiDRN6mV3owi0Q5I5u6QQkpPhd
5ThX82mBHnvlPnRqP/T20A4+Nbe+oDkM28yJtludMyhVwb76WlJJRdqfHi7ReHPV
nrjaHyBdY8fXfHD3zMpz9oNDJnLgQueUeeDS47ny3xl6gNplTJGefeCiqWjTYzvd
0Yq5F3bF8klP1dZI0W7NcymgLrLZ5JqOedFYFky+kz15KMEqt7FjVOS8Rd/Jo20v
9jOXq9D2tjoCUEA6rs5mgkQV/rWW/xA0ZKAXKfs7UbdLCbN7Q598qo1ig3rxKrTo
NbjqT5Q7tY0iFCG1lpf8WaJuntql04Q4+dhnmEoGtC4J/TKtWIiHbwo/c7OkjDc7
j9fZxPrAxprvnewkAo2MZ3AFKJrX314Qi7aiOQlNVVuTIHgaRWqzHLmop26VhtkH
jSsUdxWZSPS+6AequQK6SBQFVmZIToKGOvtAzhjPCCwnozL6HX3htGtTLqefabAk
wc9s2GnxFM4ztttOxbReIIjvErv9WDF/IDQj/WOKy7mBt5egUVNJTePuy7/+ZsLE
cLRs0GPzlvi4feiySc7jMlkQFqG5yUMaNG9VzIGKQiG79aSg6U4xfdq5Nc5RFiRs
+4ctMmZJktnY7onjapjeAGWr3+4ClZo6ELQX41RnD1CNDcxki0DJ60sURSvPXF/9
1R3Kklt7c0Q2MJ7zWVvvDgEoKhckzJBEgxB0zXt2IbOCUG+DnZCg5LYkehzoV5Gu
u4+YHuqTcPRWNLEapOh3jDs7cENQbSaseouRfQqRx1/nrT8BKrzRuXnhHlYM4Sbq
qawtCu9Y8uojBN2oW050VbWXKUirUzxlQIsuwe4OypxhNzqi2n/wVRyEKj5I7pXd
5TQAIeEziOl3t9Q/8ZL1IMiRTrydphRY3jmv9KxzYvTtO+bfW5umaEY4UWlZUbsD
K22Rv0ofbdQDB4hxkUdG8yL38sSiIXLmdNlRxBUMukHHvpqi04hnZb7cTPXMTMqN
B2UXSo9LTF7R4sYB1jCcQxTCj7e01fNGTFVik5tGDL/dLCJz3xtzqew83DRWIn+n
S0F8Gmh8/NmuZwcLXL6CSslOD/pfSk6Fob97u1CYmFladWkbBuNkWFf+Qj3XtWXK
o4jcSj4GfnAwb05XBBACMG0h9VPp55qdliLiM+fDf8Hz4PO9gu6yui8UF0zHUizD
HeXD4RkunhILdK3QJXOwzsTx4TzZMupuA5HPL8wgWPeEDe2r6hOqwqJ5qIUYGM/H
5JD9KXkA77hp3mWVoE9YDgXJ2SIpKmO2sb5owUbZO0VvoaTcCu/D+c7Nb35Ve+ok
Wx9MCzb20FutTYQPdsvTylcryq19jnY94g4ll5qeOUuAASHGe8XngwPfzqQ5SIOg
evPxq10tO4An506c4sEdVFOtr75lxEiDNYeqRqXlaGGIU4/2oex+yHnIu7HWwok6
JyuQSDrcn56taDhrbBDmRvDFBA/0KuRbpB7H0+ITXm6d9GdQMEvbeGlUGZxOe3IN
8VGj8eDzzWbK5B5bDPzaNeMtdMGNiSyKFauX4eWeZ4pNmQjPsctrdXLARYvpyDuH
Mf6/X2BYDkISj68Rux7ALgLdMBDHyaR5tI2+BjGWgntdBk7lOGswt/CF0Sk33ykz
T7peTS1zPjCTEXtdNEXlOiZQAWn8p4AiW/EqQM4Ubk9EfOWHyvREOzT2Tdln0B9W
8FFLaNI6Dou8tVd7mEoeG3+QPVNGusok5M+28mtGO28p+DtHa+dPLmmDZgpq404C
2cDZGzEN8/25sT7RlYJjX3WXvy/uXbSyVZ6CNQJjx8TLPKXVzmLuG2EY0+A3UnX4
kSjv5k0pC1BmoevekbfMYx0vWCTU9dvwAUKrAZA8SXvUj7BGj4oEDDYjN9+XgDFm
JnegibTW7QvUWo9s4IUTWR26F2aTiBLKSg1sKSD5PeVPYantlbx3qfwLtHyTGxZO
jg0etxWvOG6+UsGMdE1nj2iKs+q218u0ePlo3k4ZCspmkLWeQNPquRzIkmoYpS8y
OV2R2BTGKQbcr2IVkfr3YGoPqOR7vuPXJMJDmF3TbEIEdJm3A+uvOuBKVAWAtoQU
UyCEeXG3GtLKn1zCT5D7DTMDqGsAJ5bKbgzGzICZFdzwQBi2L5Tk7SdulaBmNV7t
EzR2EPQMBuNlkhvlK5ck+MV5bn9pa+rF1OWE1ABJEYw1HegqEWaelvhj8TBdTCvH
XbCiL4nUBVPKdCszATuTw21WVbTQK2cYEAmskxUf7a6h9UsBOLy+YL19YmQCm3pJ
W6FqPTl7lGA+V7DA5OgWN6BB9FgXeBA9c0lwQWSrYGSSVOSPIvGGq7N/eiBFBTSn
2rGe69oEJmD6B/Ayim6vE4CwfV0LooEeG4dzwsaclf5e4pBuH9ERPWUOr64ChEIo
iihdvZVnFhtoQq3yWGv+YqKQrqwuBuIgbmmbGlt85B69t79Yj+vSV2txGD2eQe4n
1HvgL2psJBM/+YJ4W3E9ZNUAgx58yUfwhl3jB0pBU67Mplh/RzR4gOdaKghYnLdM
31ggnzq+c2SM5PrvRjeTcmGeww4Xu3JQVd+aXy4J9TB5mWb+aTQ69q0H+QvaEzHZ
kLTFLzdyncrbYcrSCqMm96N9sIgoYHyXl2/GmQIeS9mqBWkwEa/j45uW0srs2Mte
N91qw9R3T9QOeD8gQmmQqR4P0a12NVRFbyNgEPcLatrpdDS0qJbeBD7llNrhbf+y
WYllGH5dAJgLWbk1RTucI6o58MjBr165jL7+TO4t5Awot9g/hK3vj2Ugm8RzR8dt
0T3MUuo8IbhbVklzlFiPrIkgSjjcVS1a0yHt/D3ewZkxoN/bGIkPC8a+2fG6CMu6
wRkfjb6NArKMUNeS6wrJwcugGqPFNiSw6R08C5I0tTMNqcwQyv6ZjsD2pT1yElDC
6Xhlquzm+ycgtYAIC3mixAy5281OvuB3na3h/UH0UT2RKKjBJch2y82SvoWcHAgG
JWpDe+7MN+d7u/8W611bISr7D9OQMWfF3GRL6XH3Nynb8TzpYkAiEqkGKReOH/T7
JxSebvj+deS9PaysH4/pCIPiNCAm/Zz3GRl+OMO79cVUd00rka+epw1Abtca0mvA
0/m4p68e/7PrLe1BwMUR9EANlD3dy16mtcXKijtp8s3f7aK4u7U5xAoCtXPt0uLE
5AE0CKS7wL1n52bkDrHnEWHjjARI0ZQU8KFJelSqsKvzb6wlCEJbhw0Ds6YPUPwp
S+GRgtAtgHlvmuyMiEA1bepBHevSEFVcWMTA/Bm0ycgRFGTu9ic8OmDgORvfbUc0
Dpx1pG7Owl4ZD4WTlh+NA8r1YABT7vAQex+tRkyhybTnTUNQLIbw90pvNTF10sHG
CzIwW6cBcxNqT4utlCGvAeCxZw8mkOgo5AKnDOqQAz2/WzFAPcij9+1B+nT9VrDC
hy00e/TawIA5URQnfsymQvbBoGi1K2FCkW/BslgKBFyFomCRgUoOdpHzL2wjdQVQ
rJ4cgKCRWkwtDy06MLNSkD7l+qQ7fJ6Qpv3n+gjGRu8rN9hbXpm7e3SO7TyNgj8z
mvAjx/sYSQJBv1viZljvaEjGs8Ti1HMAyPUwlB3hRtmqbYkjByMYFseVQz0/Aixh
exB8pJ/Z3/agSgDUiJ+p9txPM0YESqGxuyCDDeDB0qyTpydUMDCPphqrSWSuFaZr
oW67Bku8IVtTCXlmY5oaQwpHAL4oa9hTu3V9EEZjW/iSLwaaJfati66540fLDo54
1IDP70Y3w5lJMhYtxc1nc5goKmdBB4vRZKuWkebi//ww3Yol4ryn83n+tWLEed8h
aarqHSWhsoDEGSHL+fHWrF/y67L2Oypwe/7v6gj2hSdC53vCfeaXA3LmYn33HByY
jZ/bE8kkpqGJpBlmkcaum431R3jiyZr73rwq1rEFdFS2XC4g1OILtQcgCWQIwaBh
vGb8sfLLCAxKDuWyjfkbqDzXrHCrSwgKYRBsJ9zUU91UeadkIZ6kd2SYdVfCdAWA
8goPWjoo7ezH3CBjcTgl8sZ+oo1QLtToJLEbKM0U9pA2/sC8Y5IciC3Sl2wzg6gU
xNcdpRRNxihqlSbEoogH03QLI+HbbMRT0jh2vBQDWg/U4ZjUq5jjTm/DpYnYB3Uv
E2/teE/zlECEAMcHb2/x0sHRgKa8ghnRaNxJWacuniG3OVMEVOHFLPUtEZmzgYco
Zi7/iYwCSsfLa/SxEZPEsnVEI2mdZwTKDK8/XPej9uwMWKmxqSNe9P/lJzCgr3pF
GweQ4MB8tMK7wZKLAPLRorYBpkZwKEG+ECWTnacnKKpW4tnv5VwawqI6wcvuqHwH
Q5jRaWzi4o+1P6j3qq1c6qzoTDkNUjqEnwPIwtkGsOez60rW/ofZ4hIjJf5Tuy0f
q6xAFa+L/6jlDbsoeBPC7cCZIq5RxONNK5SwzmgrAZ1JT85u2qeM6hAuSE3Xx1Lg
kIkuAcK3Qsf2FQx/9v5mE8zILSu1rUITVlDqPNrTEEU/Y14WosTMqYGWDNT48gmk
Qr8RKsIhhKrLOlviTHoFNiH84hRKLW6jZQgmsETG33tcKjxq8iY9V227ZMGlxp7+
i2eCKztXQr6Zrd0QYuqPXb5Sj7zlB8cyPAR2DgO/2TFDkPJATYiDyJim5/TTa6bK
sWO9jE2QFIg2W2RchzhXys/sN+2WycDXWXbrhTIOQY9bchH7U7rRz63Bbe8CCz/U
/XVpnidqziwXRKekj57TGe2cEmqOcl6qLRLmcuCCZL9KNShpobxVKLviHZBfBdAj
oiyRgimcONmtM1p1W54n/Oz+cen2EL4paFMVA1XGH68xn6kUPQ9UY6EThUxr2WgW
m8//SUJ/XbTVa8Q7I7XC0FA403YDdIf0ga5kTkiokqdn4l6UsFJgyeFgrO/9n6P3
JUi3heRCm0dXJklc6SFmGCJYcUK2vLfhmHPrj7TasQ2Cc+0xt9vKhLULFtCrtPEF
9qcD0gN0hGiTj10+q3dBC0PTXbt2pa8MSH+aYt5K+GVk/U/FDGkHhFk/76wn70/6
k6fu4XmmxFpzt0yh+FtgmAEwG0HU316aucHOZzL1+3B6eMU6fncmjeitoKm9jN7i
D1iE+Yd0JmgDHjqtSqq9TI67wG1RjVwH+KTih7ASJbvZolw80i+1gZiaPniTd+3k
vtVWwOVUi/v+ywnJK6u7qYHEPPPFtX/zSB15EWpw+x+jdDgk1WoLyAPtZ2FogcUv
5u/9sBCTvWnYY5ZeCPd5LETMJkiNpl2SJ53vbQID7udmOyfW0l+hcrPVUGACZ6P8
wf+7ArzrecrZLeaEmVmDqTIOw7OMByBJZWb34ul7+YixD7PjhnMnF9UXP5iC9kJP
CWUFbEMh39c4ILTnw3hgBguewC04lwc0O96rDLU6di6r8as6Nw+77bb+OJ2wzhkg
iQ8jd3Nic9UX9T13CErUFgAXbM2bOBx6MfiW5VwicleYZSuyttsJOE85rR2GGsZo
XUmOndD/y6F7jfnuvFP8SuxbxwJTGaiEWLGzZ02tGErhU1GbJkwCdjkUcw3WbTlu
jyBK307gcNFaB2hef97TtfCFj+mAFViH1prQTrhGP9ytPSo55g9lAYKxoA5n6wsy
pRmrBuL/16ICuETrToU6ECHt3qfFXvOLRdEnAVpFh8wya0kvveuMDwErYuYa/3Jg
iK8vxAk/vFTdt+EW5Qfe4htYq04Fe7UvN7pgwKN/Y2jtl1eBkkUhEAIIgp8t7oOI
+zfHfHw0mCVa72HShVKR1SZHP1gsL0ycwo/eRn/CsrbTl2bz+CfL6yKCSK82DRTL
3SzzTeZ26mzHOZwLh/iY+tZ0bWceJx98GskVL1V71aJprC1EzOIAxhEZWxtzYiUC
Ko79OJrqCgk1qd08GUvGcUIpj9BisHGShhdUELSlLg94Uu03kUuarmI12HLP7ctE
2LDKqtRRtScgDu9Os7HKmM0liNY1SXN1r5S7mvDvZKyyjzf4hnEAEgjrhBQEDkOP
0FURXL6U7DVI6Whg5tomY2oF6SPR7hqbF8TtCZ0gSyYhCV8hSVUCr6swmD//Cxvy
8Nx0Zqc3f7UZqazY31Fx9QBFy+pQC+pkegzbtVhWkWSofKh/5ECAoVEdwYpgeTjX
XIJrJ0bRaL85cccP0C0FU89d3ZqbJzTEDkhtebGw08/XB1wpcSd8DHx0s3p2PM67
r8OXvNwlJ9ruf/NE7AR5rzATnb+LNY6guWVWnJXagFjI27grlksfhA3W6lBDyX7F
7hElyt7+zQyiOL/yH/n7JP7RNIxojIMeVWGWYpX8knuZuhjMO2Ytm35UR9iFYIN7
ECLFAgcdLbEJvistUL49UfA1tOYUgG3fsXStdQiac1ZgcrpgA2U49B6ZwjM1Q/4P
41kFyLptMjMHQHDN5aYVp8CzA0yJm8diUTh9+oWxOnRRmtJcxwnoHRlYYv+k612I
EB2z2DywYsCX50tQe5XYOzE39UdM+tTiL3UvFB1jOH7MyqpZ3zjurhlErNfpBz7/
AjD1IFWICSo199DOYJpzr5MJmsqFecgpdTfA5rj+NM7Cp9AvylEvg/Q9qXQOpFpJ
OXu/zevEsKju0OmzpWsWMMoshEziv/oBYsUtxS5oVYXlvGGw1xJMDqqsWQovV9uG
Fa+Ohy+BDY/2PLFhXmU+Jt+5KHLPo7zLBIoyx5MSmA7Cng6cbGdjOyMjIPWnJNtp
nFIR+eZyhAxpE58kn/FokNIvRIjCBd+SPTkmwhDUdyIndzaWwN42o20MT/0f/NDW
rZIqmyLFEMR9jSquYA0EIDaKmYz8pveselWAiTwY7aZUMiQQp73+ofKUbOTNUmzg
FKZ76HwnB3JK9LJh97TJT2K+UTb+jizEgvMHUcFeVqmWOEBg/wBqHMGeNkkURAjZ
duCSY6I1DgI/hIl6ARLIWQ5CV/Vy99DliKnpkKsAxMoYa1a+LTIQY7TVwj8FWtG2
xdkJvg/yQ7i1aqm2f8dA3fB8WQqz1siZA6XN5KzfTaAC2GFBQ8KdUAtLJv2/E/gL
EpImz1titMXuOSRxyUYOi2q+7UzkSKzSSbyg7rEjzv8/RNMPdGr0OGfLHaWm06Mq
CDBW6LvZGk8VRdlkkVyL7TKdGb3gBZPilKEvZi1800orx2nKdxkmrfwZ4ps7lHxj
9GdqowS/s0bh2Zy2qPVKY9tPR5KNIlTJRmivkM/zcEhlh2i54CO5H1/efJzpw565
N0QCzHQLL0nDuIBt+hp+PwuDmyNH3t5TkAHKXtCafvASQOy2JeHLI7gPYYbHJypn
gFq3GfxhRsKqfP8nyHvbzZc5X1k6l8qDT25lBkVaMtVsCUD3iQadcdEPTdpzr+fG
H4hSOOPgFih0TLppBeOQeHNRPfBI211cRctoEoTEDccd6Q8kdmpFkVg2rukyHYtv
Bfdq9Zngxj1j/5ZqhKxRUMxfvt1VOaOciKdJaveVT3sd87ggbbZ3i+FJmKC57tJM
MKVr/fX7Oa8yDK8YwpFQ0h7XmSomP8JbXUR5d6cZWiqfGWC1v9w7wMYusry60b8t
mdT4H7mGvJl3DaxPfvy73cVs38o2S2jEyYgJkKiplfiEyuILURIMRYNZTZYD3WVj
GXMirp+KlNp3DpcOceHzLFwga6kQPk38AztqeqAHVsJDe0AzD0fMqMYs1ex8ZxWP
e9CH2AIaupl6WzhJHf5ydhOT/ZrCYe9LG4mMg6oYtO7I+3vaguzNuh4duVq365XH
1Tqsxwp1yhw+dFYwkTbifOMEXVsrjB6H4ZxG80ZnHj80drglSXwMULSGO9cnEXOl
4SltPnyJsCmnnAuiylaMj+MnsyBjRH4fCqORNaEw6iXPqbkSBQHBIq03YBlSazJT
5WKkvghma6FdIZ+CcnaUr5LKOKMb6795Ln5DeGUVU4IuTG6l96vHoVh/YDUVtcld
2qX+w4XW3ocEw3WxvHc08Sr6wRDbN591NFEmXJTkEY9jYaBIz1OPUnu+GMxWaKCx
7Yj4VeLj1v8VaPK08lcX66Uv9J3pglvNuSQfYDv1+cBAzwT5Upn3LLJ7fE2Fbr39
BCd8yNO2F3AMY8UNZd1bWmiR0QWozjUwXIAn2f6dzvp1IFmAecqVa8ZysXKicpIc
NdRbNJFjpGRqpGBFfX7+8tvzbpkwM0qBtwiTMkbQshNnr57VjSFA5GpHRYSdy1/Y
FGgTeUIy2HV5qIeTYWPgNJE+KZ5gFk6zGASfmNOHwvJRVLMD6UV85q5oaXQtXWt9
JDGVZn97rS2yQ4141AX7R9JBvhl9ZUInrxO8bu/niuMr5SatvvA3p3aSJOn3xo42
4XiOUUoP9wYA3ZAUsHQzm4Ue7f2Vpxp8f1FJDbBDT8cy5UBw1xn1q2g25PMXpqKh
XvTK/6oOAziCFu2NpXoOAkW3a/ON6K75y5aDpjKsJPV9eRnRDumT6i8w0j9eDsjx
O8tQoQC/YB0X6LkVNY8cu/vBBHgA9vUdzIvK8X8BAvYPmzd/kIRAritbvHxx91ez
p0Mzhi4ytNPwr7xl0mIyEAfHGZF9VZKxnRl/lpR0E2zvp9QtEjis2L1FmCNmpnXY
jcRo0nARGEQjpnaqwSROSfTEtzlCz5gzr9dIxwr75CuVXYi7jC0fwKmWyx9UtZqL
miCswo3cG92lD4iJ/D57MYarLoNJddcguNq44KOmvqSpEvTkOMZ3aS3mTqvepEj/
5lY5a1vZ4q52F0tCUzSAeyXe5VXT5JzKsq/pPkDUdX4nkDFfwmWnucGpp/gifzuT
K3ABaDI/rO61UqS0ZvZeh3B2xQTpdHYw3S+7lKrEs9XkAtfdTqVhUalahN7JcZEs
CBsT6uQTzrKBXX5Juc2RDhPvuctNBUic28siq09O8w4MVcqmJJz6wqCvChxRMxbw
s63r/Kh5ooGUUJX70DIfQc7g+PfvD0913AlVBhk5GcpCavTzkAbf5iVwbhbrEmT3
Cvj5ry+doVxZDOFFetfk6+EJD8U7wPXK1wQ80yLqLS8iOwkKFzVMXmvYIQGp/19F
TZ8fEvbfvhAu0hCGi+ielUL6o38te+LFF1TpS5n64IqkcXdaHv/B33cD1Yp6UgsP
v5k7N/Eh5WW7uyntGscLLT/DibEj1NqF6eSOM6qAlumFkDrfrKwlAqu8Lgf9g0QM
D56OM5wcKcIvvBI7iAb0G3Cw2ueFoGZeo9TEI4nRtdvZxgmqQ4mwXgLu+lUGxhE2
bmHU7OYcBRJKHHqtdvHq7qsPLi/r7ZuhLOiEhCDCqnCBvElTaj6avCPgMPLz6zy4
PwG88j1tUi1xhPeGvCcGk25jxjRzKASbj8ZI4RUkycxBbZitzTq4Jpp8+xns5WQS
KKiL5J/5X4E+8u4a9HCLKU1U1XBPWbi/xJU0JhfxDszijYrAZHk4mPmez4HXa0EI
96ZCW2wWhSTwdc+11TNcxf0+k0GPqLVZ5SxVN+/OuAMxKg4/iCLYEehZnlWcFpr2
IKM2sOsfeFt8/p1DTMqSDnKDz6HZ8/pbtLECSuzHr8+iEds+pafy1u6pFcbgpLDW
oeCls7pEyi0CBDNnhcGgilRgKz5mbbGxZ4XuAUQXYHDgGBIn3pAKo6IA8Or1SCuD
Bm8n58ucog+lFinXnyU3xO0VwJnhACwLclb2/4w8KQMJJLze5tNiupq5oB5bEUNN
dOe+oj1eKBmvg6JPvK7N6omvoLBSM3P+I3MpTI+Pf/0FbF3TLLdV053oDfpxYoI+
LV8kkAZxrSXFeP8wfMG5js06OvU/mml+lA6BsExZYicpC9CfPm+ATG+PFNbz7o3T
eVr7LJQh09/d774zrlYLGLYjJP3ko+iRYTLCRC3e5p9I+HO7NFBvKOMImUFSx7Lx
FMYrci6k4r/52TEPUhB/ndRGpRicbIJ7NHPfbRDMXQC+uE+2jAmj+91LLE/tTN++
q1i+by0haghKz6mlWW9w9evkDBUbQ08V5JD92q+1gRb2TvPOrPulDl48cC3IDUqA
oGp+T3CMJp5Qh9Z5tkJ/MXSdPBeqLVplCRbJCfOB7PL/y3O7+Qoa1P1MIz+Hpsih
0LcQi4ACVLj/NXzjfXDINeuOsJvdxAxbPxxHpetJO4t2c+wgN5zLoNqrhLm1WAAA
rMjeUfeN5j1vBXJdr7LctJynTMC7CCHtV8g3Xm8SI8pFYCkbwCCHzCelyerO1nYg
gxbTEow9UXDOD20cLEe4B+z4wAgwubGsKSwNFdIV3rLXWfSm9M6u+Z5VxfreMuMv
XY34wjDNPyhGoiCuzNRyhQG/l0Vej+SjAPmUBLfMPocA7iFRJpSDO4UHt0PLMBgP
zgvj/WRpbq8JRxXUpE+u6EMr1iTzK33RiV6i7bb3RhOuP3RvfWzSRgWA/pWbPt9A
8QTjCRp+mRgrvixnfYtphCZ4oVfLoNhjErPxuGvAmWFv3vYR66WdXJ78PZCJUT/K
4ZaR23EBUbI1DDuQVH/AvnhNhMKojHNoY9eNazLK9mhzUHBBJmlPVza0x2mWaGVY
iG1iiAZXqz/QSC1U/gL44Er4ZvXIFYBuFW9iU6+RORdf2rsCfFLF4g9KEN7IwPyZ
38/GXVTTf3HxVRwPqRKbqa9+ETCQ/+4KcianxBEurkF6lv39PX2pKIyRsauhgRkC
CrRQUeAseLZnwtvYjDrkG6j4qkMGR3ZG1LUG5DZDuo82MwCg4ogRhm4aGEXI1LJ5
/FnrHV9BR7bHJzw1zabvnw2mJN78b+/mST3DkfCpy9dRR3W/l/tq2GO8+wns0Jxx
DEqnCac3CFXQZCH0oWwKe1YA9R5z2KtpstSXRc04dYTv/lOygKWa3qQKJLEUxKWV
jRa6dUY4ZsbZHFrH+Nxmysc2tm5hFb2Who+YjKn/ykrqfhS8q0luQnNaXZ2gETN1
jErLsMfPFGCEyHX26ONsASGpI9bDWmFILTVNEUjlidM6olALgBxy+hHiIrMC76OR
zrMEacUFQic14Vyyz9RS884JAVILjt5WKW0iHCImHcLY01RF6upMzvn9OkAm1K5Q
mEFecENIuTkQ9l1qnEOanH6bEmHRopyDyS1CqmUeSuRTG2xsKnr41IDDihKBYq6K
sVbPC/HOQ+70NLeZiUowyTxXUn5SPaJh9srGgsQlB+2/e66uAyW/L7+FEvIQs9lK
vbpftuPbDtDeYirl+5gJywlWq6p4P4gDlUOUowk6PMeKvrs0j5aCQisMfzGsCNhD
gb7fDftVvYhc/PVWG7qiR5U5M2eSzkNalHOcbqH35oqPh0fRkciOLbpnHql8IWxa
QNpnIXMK0mDoX9LSIJayOBJHJ2J547ukp7gHuulaex54pUjyVR0s+oy2TdGIIoY7
YXg1Ge5om/bM0x5N2QCMd9EKEcy+yyBXYr/s4zYF3Jce+TuLN9CjGqS3yLyFHSF+
zxRtwUZyTZU6bkX8O/B/Ey0gFhVKZ0OkM6j/MkkgqmOw6YCDaqJZaei5xGnIvg8D
kIteo7jhcXWP1HE6hDK6By71A4j2KRBq4Kf+enbSEtVEWQEg78baMYyDSzs/TmtT
zm6NoCVuOyVPHcI4DfhoFY9NziOkNg/l0EVXhiTu7wsCBIcb23eslIMMJofw5fyb
Y2cgu1TO2bLKGRjVuEyTEKv17D30EfS+rQxXM0YQTYvx9Ru7Cv2iEw5skskPMyJI
yt1CnyC3tr18sIuXCsHfQyxZnrp27o7wEBbKTO09/+EcviLBuQUDdUj0mKFxSaDj
Trz+pYaogQoZjytvjtd3Yr2P5TSEpCoZlc6KOafcCGt0s+cM22js3mEbF9yJsZlq
Om0xLPAwpNO7md5aE471NlLzcIC2b9+x3OD9QgJWkvOmd2y7WYsU7znQbQOGNvLD
EpqrhP5ky7P98kvdlXQBrcmGyty9SZlrJovLIm39sVK6eaTOob7PhK1E1O9iKrU8
qUzNATBM/o5fRUksNSYVt4k25wf4vAg24zYhAQfWOpUp5suIRydYUP0f1fSDyDle
MeXqXL9vhtCqQPBuT1si+r9ZnH99sc5WmWgSaOq2AUeQZIhZgJ19XBikx1ICEjyz
vGP+s2zUEbfifgVghh6BGfFOGMuQQ2woVkS1iIlVsiDkAYQGBh0VNA/xAW3hWCHR
bOsBr19BqEXGZEtx8R62HPreq3HvLDOFzubWdbGV0ZsF9W9maxDWsvs/8V24v8bx
q0LNwZQApvdWXtD2tInXuNOEfKt56cNzU8fnZBs10WVYYmI58OqZPzsJ7UanxAVs
ssX9S1h5j+ewjUnKfbLXHJolGNO2v7btwJ/1mP0GOc6/Ep/MDOXoRGt26IHqoWCo
ZAZmDH2AdvUgIy/NKekQxAVyRrzY8JtGdpHVFmYEJLnHbYCel+k5bLPI6d4ZFBWZ
TpPmSlj7UDMt5hcv0dJ9i6rCCv8FFMyHsNmySlyvIPEhOZLZ9rqKbG1cu23iB/LQ
ureC+dqxzvAWoyHd2oqZUOqF4pb6uxaVOlfQ9W5ovuYKcXXafIqcKx++tptANoq/
SGjydWzvcWcokUMznXedJVjKT9g+bt40M6NpqraUCoGgtwWjom5DHFGcCL/WsDYi
KYxd4ewUpqE9XdA1k9RIHCR8K7sb5tSX8V0KnUVmVNv6seXCRJV8syumZN2m86L2
h5b2YR8lGC8+hla3kGiqlgTfz/0OMFt3/x/+ubYm4sPplDVo66MvdmI9jsQ4eWls
iYTprRnriMit8IDEzqM8GBSnW23uRZJ8FjcUkly3wNncNvgaZ7B9BhguQ8txBEi5
7Cb9ZRiF6sdkpBQkGiMTojdH2vecn/ydmNEx9OAeCdBiIttGWuNh+hy+WRFXiZ7A
GYEwB1TV0x0IAVn554Lp6fWnFLyOmQpOPwHzaxHV+p3zMi0YXR9X2jEdJ7JZGTHl
cIQks3sFDULinEP15KUIVz12h9iguTL3nutrpfOhedVgPgcyjzKkcqEBRuYzSr5e
TjPEkHjlvk18+kjt5DdyqDyfMtLNt5PW4GacHua+qjpjDpwtlY24jbr/6h4iYzg+
uhV+b2fXJIzNcfqBC/qwu4y4YSzHW9f+FYakBd3r0Unff9HUu2x+Kn48UWlS2p/R
7K4QhGuwwPXaalqIUPLAmBbhkXkZRoXaYv3p/8amxQ3YnaCSk3l4t0GjHAxLa/5J
SbAuiAjarKrlLRwtHUvIec7y9W5gkhzo6mYAXGszmV5h6ZRt/oTpvFl5AhJij/rG
Wy9Wy3zbz9oHfw1ey6+E3ulfrGMOSuVS6/9+k6T2FB1zBkSNdY7C0hb7EXSubV2K
S7GiOLQMHvZFwy5X6yD66WbAkQECzHhONlDP86GwkT/KVG2Vumll+fswDo3eN0rQ
OBAa9inGPNrc0a4YwxyIBMjIa27lCQQZLXEW0gn8YDQOEKwiCvPvAuY5BqgLNn8N
k/EEr6BmX6BbYE/hIjgiHCvxe08huY+mn2kd3mXP1Lp/ehE5mkIEkpiZyqa1/8Zz
X/phZKMKAM8hJixKCllyIWY34DDn0P/+iayegglmd+7F+vF3fv5cjiE9i7QgIIMz
e/nYMleihGqoUHah/Evvq55OVKpNcyoeeP84f8p15k+8M+pJyQjHFcozpSn5RXSY
5lq3N2SgBeYs8MrwwBi7AwFenxL5EZFLGbZesvpiLckPHsiMTeOs5DYUdcUlmJ74
BTOTCLs+A/Qs+UGkjCWlPQ==
`protect end_protected
