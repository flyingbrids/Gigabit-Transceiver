`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
HSTLPtDNj3JKUcaJ2dZRa/1NYv4Sk02AJ3uSM4y6tcnsHUDF+AE7F6+9t/GSHQGX
zm57/cYDQ1Krsit1gFCzJTJFqUevfQi4FQaLm/hx//4WwyxBOdr4wjyMJXRh4p1P
Vgao6ZvcJnidAdzuFFUQQ6/vytWsl3RXwZzWnXpEH0dSm19DyeAhcNfwXv7vj06/
tzCIxDtmJGcAD/wUU01W/+8hIgFc8SKKVG+Wv4SyKbimqImST6CnHuzeoOcUQcDh
pVGoEwa7tMow9bgTCkw6nmiztukHGthCV5jPu7KF4u+7ir+pHH/2QF830+2XblzF
n5wfeLHnzZdQDGbtPeS59A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Swb05jpmGeEZY6/Oe6LO7cZh0F0+3e1eJBUcy6k39Hr5hQCGO47kUUR82MnDIReT
yIpzTPuScbx/oQQjkq3YWH0Vf0/Vdzix9wImh8HEKJJqxaccAqtujH0ZblWyEQ5E
IAOdUPubV5ouLbjvawcRL49CRjf40y9uV6gmlKF7lls=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 28512 )
`protect data_block
YHd2PpXhGPHtZNaaDumfeD0xsIpAW6c3+Ox2yEGUgexeSATluKdpYkYF14xVch3m
aa2CFOcdL2maqVeZ7oX7h7FDd8ax05gses12KF1R/oREUgfModFlH8tRJPqQXzQx
7mv855f1fvxjdIIqnT4+gUyBtfKGUxohwSDTL9O/aaIYyiw3PCx2Ik9dqadD4XFs
TQzKXkGhBgleeyxRl9y8jy51xZ6iSUyDUC4W8Afcf+qjee3KC9pK1T7iHSCT6oCl
dGvIEeIW3JmaAEL2QLMoHUdiabMfFMTe+YilO1HHEehwwT4MMr55vLK4qztor2PG
YgF2PGttfnIRTJRth7iDb7iL0RuSv7GcqPYQ5Y+N5r7Inme+8FE+iQRA6l335YoL
MAoR1QnJHqyvwbRcRlNPFTvHF6rjwmg9c1MLJS39Dbci2Y7Z8acCzPC9eJGJrPCJ
0206UPA4uvR4gXP2sUbmuzSouZnx+q9WLIFgLhaiwt4OSAQDiqRTGeevDO+wvz5v
euOLYVK/2ON6ABkZTPm5yPn8L/ZMFd9X2I2eEqvo9257/mXQIyFGwYfQIe2Pc2IZ
f3IjRgcXCpngKtYRgA6+32we61vD+czQN3HAKGxklgVBsn6Y4etlsy4w16CWpYH9
28t70qWkZ6FEFIjq6Ovf5FzNBVhR6/LhhRZQkoMI1B9+cP8QDhJ5Gylur4WenJJd
f0Cwq1bxUXTLIVOTUMM5G2YYnX5JMOk+enWmFY7v6fuLJ1jBbbzHgbNSlddGEiGQ
ZGhOTg/1Y2JkgyIg8VPVLvGKfZkhP15rM35dkM/EPGftIwEx9WNsbtfsnsZ6Z16e
iFTCSr+tvpZjqiMlF8XSgGeLtCiaJvgp3syPsBARco5V9jaVjEnmWOmKEGaIvWzn
tQtCXfdSqk7J/iW+Tcm5V2YxSBa4ngD2G9b+AZ2d0r1XXA1zgqS/R0nXZRdEtp83
M3Rm6CYenmkgk8ha+cEy7AIVNfi+HkV2i7w4y0GrLvXVIh5g67IBWTm2RPRESl1b
d8K7rENYPk1yvP5blEr0Wl7w12I9XFEHPfr9q96yrspvk8hQT9lvzgFFNqKae7oQ
EATttrwgcH5EwiXgyLRjTRM7x5Y9ffrOjuFp6TWx6dizZiPY4BiT1RHS1ybfQQWp
Ctsr7oDUiGIihOkzEu3zUbk1LHtS9FVYoGBnJtcnGnN1xdqcdZ3P48nsUQ3zzQxb
o9Q76Kn3Kj8+hYRMHYRlw2MvAYF2mvjMNyXlMWfwIgaV2Q17vpA1mIv24WRI6Xdo
rkdb2/7bXsK7XHpLj8ZsKaqWrEqQn+YJSfuV23ynGz7HSeR++XvKiCWY5Oezs5ko
IHO3vyJYc484k6GllZGjzMsxi/MwOu3pyg3rzYkbruZYP4xKeO71io3XrATXfknL
WciTv3+0Cz39R2btbDEKv4cBA8vC2h+Kc1//qHfx5PyFuhNEBIFItwuX6qx211PM
C0stb/znwFkDLMC/Zp5n0c+QcaqpUKQ0McO3491hSjdDo8Yo19v3YvfTtFuvwciA
IUofwUCU3x/p+94McJ8cGajOQSM3kFXB1FMl+XXrR8uGVcpasT1dqpJ3zxfSJKPd
WNu4jFISVbLpPpk1HkVbU8nodG4SHaJszVzDDWvvZSBhm6kT7Hrdm0obdWj3Z53r
AwGG7XU4wccX+bDKrLr0nsLey8OHZmMVEs5H/9WpPFDgUp9UEBFxVWErMe1BEUKP
xk42FkvCfpCXw8GIxFAW1Okf4w1+8jfGGX9mazahKPwIBjeXVXcbEdrTEshFgq4+
+nxXIehtIYyR+qrrUMopeofD7sedwdEi8pwoKmHUE/Gy/zMh9zChcx+vyr/7hbih
5bhaTw20jiyA88ZHmRg4F2AfVCSi2SUoBa3rUfui7M7NuX+wc7EESOfjioSk0qNU
UvM3tMeF+3xo5QsJ8G2mhfL6EAI8jJA2wfYTn1aGDxlk2NSif1IW/IBZSbOTa+bn
/s+ky6XUDeQPdIhl11rgV5+19ryUVS2t09gvnhr2hVm2FUPk6UXQ7VooFm/2Jc0i
27m+/N8b4MsujmpFtLvH+n0hy7kF7kyK0t5MTXuS3M2CEKGcub+ilnB9ep22MJCB
h6a4u9ndmbd7/Wa0CB1STMzFN8S+Rzu/yrGZbQ5b/90sIHzaMb7k6v1QgD8wJEdm
WUAoLgisftqb/IOwWXZ7Mj9337d6PLLyTsEGgh7ChfWbD06b2EQD6VSfZ9sMi+6N
igGBB7hWYOoHi+WkH4o2b7VptPwcneYMPnGP8r66WyTDsjL6Rf549Xah0kkZPyeR
212jlLA05CafmIwbtxHEPr7eNLZFA+FcHcKGa2/98w5o9MCGFzP1E9XKoMfXxaT6
a8sJShShZPWiA4YbVSL8OFssLXc8XbCiTFhDC8gkU2/H9F3hXxcfQKRhQnE9QV1N
59/K9h16x9/yNSKpNX57CKQ4xTkj9cfp1MQV9wp9euFWI3V68reA/SDhkr/7GGhj
HvuDKSPA/nZOmF0xzqce0QZdrGxCSOK/uA3YPRxekWaq48VG1gxrwkhplwNRoqaL
a7PdZQyHYyExkpyWTSw1XxKjn+nGDgPOwlJvIB/SFMr+iH8QKCoEC1K7bvoRlib+
u3sssrS+ma/hOeQ01qkRvcs3dPpn8HGxV69+/r0bybNtRwV6DiHNgerouRtHbb68
ymAoAfhF4H6afeog55RuVhFjwslqmpvlClwu2HorIHnFKnFB7w6G19qGzoT56sMY
BNntxd/JEFbQUOhZrAVUlVibdAMPNYxa0ba6DdWeNE++Ntz/jJjqUdGLMLtJwNAq
fUXs43Czi7Cu2kWvZT9nFhVKEyZVrdP5+UEJSTaNHeBIwG3Qgf11ml0xwHWvV2QH
yu4Wh9OGox7To5Bn1F81GHiMGPTTgy0UZLVrGXYU8VufeUzVCu1Ydrr2jBOaUdw2
/cN2b5LGjrDZ49iB7LZTIzlXwuC8K2C8i90JqBz4QTrQFahEXRQmMAERLDrMKw4j
HPNb6gRh5oLbolegSRXZOldPTREdO/1XjT8T7ls6ADPEVYyNLKyXI0A2+shKoB0K
R23+V/XW8x9moYLUhJ+LB7T+GmNHcgcHIDHapfEFf+R5IlnXidgKxiEPizpXT6Dd
tk0Voe+I/hSv8kI/vJf9wY8jty2V9zDtqhcflNH8jsX+aNmWKnspcY5wT69JmBxS
zGQ2roOiVwRARgEhFD8sF2qaKiFu1X2m1bmOtmQRIeWb9wrJ0WBf1PDbzjer7FVG
1VYx6QYNeBSVHkWQEqHNDf2UtrSmbXI19HH2uVMr0gQgblNWyTD2d6ulbURehVQY
ye6mfN03O3JeZp8vHafhnZ/NLdLeB8FmfutRxS+KVPSy6Edpg+yL/7pU6tV8bwHV
/6uwKlWUjBFrv694ZTRhx83v4B6v5UEM7t2AhPRbNeQc8MXctOqQ860OxKwVLann
O3dZL4RBu+qkgFQZjSBmJQPLWNjdBy1qK/6H9hQT2ncb+n21bPY3JgxsyL6aqfHv
FbJwkABApjdyzkU+5zRZIWsOIewQO8VGXxN8tgakA9bDNd3rwIk+/SwYOKpgewvS
1e+BhE6lti6Rr1mqhTRU1V2V25w0eqfdfxPPBa8jUrnwEBLZrJkgnSiOb0RFx7na
/I4OCl6qTDR2hDUnt2r/hU3Qny/wGFGyM1ft3CoU/bbJL7yNDpGFT/qRgfhAyMfi
A/KF36TucNPJ6vLjTR6cCjbq2Tqplwyf6yXsTA/SG3sbp1UP2g/C4BM9CFjzKV+o
KTblpZsImeyCSRgB3vVG3M5jxMwGsQO/Jnf98zjNj41CIa65wlFckz7RCkaPm1Mb
KcIYjKOaIaDmbRAB9FvWYvABsKRd7JooHjghwBlIrW+HUSvCQnkJHLB7JvDEvPBc
FljjCkfjQLbXG4Sk/O3uqxXSRDR9m8MjXmw5oKtKSZj16zAAA1tSaAbIbWYkFSbn
boxY3GUFl3nfisCJkcBKCsVsAeRAc2TuGXZmv92EZCnxHJFJLSr7fl3rlqYXDLWd
uTJLAwbZytFMgz1XnfLzn3cqxNBRyDa0LHAMwdGca8MCsm95kiDNM+d29klwQspA
Om1pqw0kqabLCPAfxUVo9LDa/msUfwycXDDHD4AK5dyDtbSNBRr4pq28BqAitcqt
Zt7bw41Ozfx3zft60anlLDh2O21fD6UeUfME7tItW5OBTQRPN8Y5uWVbJirZgI2I
QHKl4hvQVIsFujEag+lOIvdK9jAt9IwqcipEEFjs3rkpvyl0YkGbUBIwINAl8Usg
77oWUBixNJXKN8G8on5LGBifjNN0efHhSlJt01sisza3scewsbEQUPe9hbhByn/V
7EZg0uPmL3okRG9J550bYtjQm5bBXa1ogqluthqK7fdeJDEI2/tI+e96ESk6F2Qu
ngH5NXWuvqZGnya/JAwoveyGIvOfjjMhBqFhaLv5V2j6v5iIVPgCq5kznuzrkUUp
mLLrkdRFSChMpnX9kQ8stV5VbKuUGQkSBS7iWMegRKb1Lr60fp2hjes96s6Qyuli
8XmZm6dwLGSFtsNNlpE1b5XSJRyNHeW5uvZTQeunS+FT8CPh7zjUnCIU27VjLzyI
pakuTtgeYxLhvqSRZifkzE49lgdIid7FUU806k1H9ykXKoWpBSAXGszYsrahGA2i
a/1q+v/BL/DJW9lI1De+0rL2B8dYeblBjr3KxPJg2P3I+buT7nHn8KSawPYxIed7
B8q2mfhD7sMJ5u4kXNgnjByeTMbQLCUmRU+63MtmbYzSsnE4DIExm0qXmVQj10yW
tpfjcQb1FoihmTokJvDM5+I7yLLX9u94nN+o2s51h/Z8Yr+XEqycTKc1OK4+OCfz
NhPLcBXgH1tOkiOWrkqfUO4SSQVS80sAMQbIS28o85k+fFSPn9JBr1hsL+EMYcie
D8pi9f10BWf3a7sirocBO6rp3N9h4zberJPriUQXokxG6PCuECmYKfCj5Z2Wwmsv
GYdY3Mc8FH9YsnwrfxdOjYGqHankcv6yCtVjrs5iQHJb/xs85/Cxz62zzMNJo0+g
E6rOB8gmHEJXCK9ZqY8Mmbid7oZvRCaWbPZJWX4gRyPJ84dTABhJsyzyj0QN0P0s
R0HzWUpMG218KpYhbqcooN8kWlCU0I2y75sp5BpUgcvOhjvYmUQAqiaKzHAW8zNK
PkINw0H1W1TWGL4KCZpNFZsaTYmuZZpOxf+srfYHt4bMlNHc1ZtrNo/p6OmXCpdW
+IGNcqYPe+fO+3VqFyUhZk2Nb6P+wI9d3+FNk2AevYhqugqQn/due+IdsBSjKd/E
rIsN3mpTjH+4XYehkVpiIbGNiFORwAe2TC55xvv80PlRYsuXuOG0sgViPNWd8Qle
WrLIVnwQWaCuxhfvQIf6CkWw9kDBDnlbqy0NCfXSRVNyHtwqZYeL8xDORbjZC9BW
MlovjexeTyENrzuxUENNUaLHJuNdFc04XgK3ZBVoyBYedqH0QHeJwZ1WjA3nQVwb
6RIbgEL6XPowkBCLs+0Mpg1dmHB1HWLXGMx/Dw1kqN8zt5uAKuERvMRMTTklghVk
2EfLpstavMAPy18K//gSOfvJIMsMjzcr4c1lDGXGCZVceurXmabAaZZocAuobgiR
aoq2G5t2vRKifRGDPHfNgtyh9+UBCK/BIUYG//239hHXu9/0Xcj+M9Xd+FjG0Chi
r6JsFIGuJdtKasgbUGs77okMu07sC4GAeet33jKqXDMyPwXt4OKUVt2zivposZsX
x8VMaLUYRQXTUFqGmbtFeauH5zQBdkWMX4re02zsZr8D1KWCVMc03587yfvlq27W
OWDzaW4q3RCGm3P6hoq5oT9Laf+TsgCI7mgsx7ZzNVKg7gZ67uUkPr4EiMqh/+Pg
C5xZQc8l84z6c/9qKXNsKB1ff5ZaFBKpaRfryEOL4TyfNn2C6zz39tqN1MFNV36v
Rbw5Zz1kzzwwJEY+dyK41b+VD+7XB26ZICZCvsXwL7pwhTmlu5uV6G7lBQ0/J3a5
gZ9LeJrvEeE9bhMzjHZPh7r19mC7puP76Gjhs/vKFoASk7fxLBiSiruObIpvl8VR
xzT2PF0ubd+DhlRjS2QgEehO966D4D+LK2FJUoidmeyMjXHXBF5oKnwuSHRT71hk
NdbnKIvvwtz/9dVW3oDG2DaAtVFq8eKHVr5B/LG7uSMassbl/FJ+nraW2MCz/cWL
wlbM+Tw0lZsnRF+89qjZRInxzoZKuRkpWhJ8vdEouXMseqbImfKseFgTlIeCbtII
V75Jm7tYbnAUrSneQhwLfmDY6RD1+J+Pu6xIlRw57uKkgIQkozPYNrQd+UrQa5qC
c7JA1uJXV0eoxKtoF2ts67sPAykkw0xLbjOHIXcXddyoNMGGg6777+ZYf9xKMxwN
yByOjGiOTHXiR2eQYYjqowl9bqdOpXTjh3R1Gm6NwVvQdtHbvOuvJNOVjgoXBBw3
BDzd70JZoUBITjnCVN+oWsyJ5GyqEHerScSr4qfaJRB7n8FVAa89V89JLUFKRsiM
ZD8SDw3yDosZZVRKTs8bga+S6fHPtLNNKa9qaEZv0iNcJxzqXm/pFOsF7tNK/O/W
XG3FYbwzfKoBXMK957Xg8gAitwKEka1YwYUBsj60vchFmoVcU585O5/x0bjyN+0O
vPSTQ27Ki/X09bTRe6VXRzcHbO4CI01xT7EmcUIEP6tOhbDfeZfDmBkITwc4zv0v
7Cqf1KNTmVUbhVhRP314FjGxfE1DT24rhczU3/oeGZYO92392EOqBtH1MivasbVA
N0GH72XxNl6ct1ZMYQX8Fwjcb/0Cg1bG1iBAPARE8v7ss3WtN/r2t48rbq67iaoj
3nqLOdRaGV8l99O4PXYu1IBuxanxJQxTQcOHn9tP+riT6v4HOF0FLQONTZbaNAq6
8v/eB35Ns4RV8yOqp4L+eznPqg8gpjMnHYAfCfcMLc8lRrOaOFtN02wKPUwp4oig
Vyou/4RgjzmClUScXyR6tGiyfIH1f3xkAqLdNsoAsgvfZblMORyG21YLeYfTzuks
Zohv/VGsGHRFqwXW2YOQxg2Axk1ethbHYszSnF/N+F59lcZTFn3nxM+nAS19ej6M
5ehyI4IK08hgiCZqhzVIqbhdOrH6sArkHHL/jBYSWck2vDgvHqJuVVh9zsQ6rsiS
cqodRZbrpeiOxwZJqdFFL9XDDYR/b9eRQm2ulOTsKdDge85vEj8oblRPhAWWS0pT
JyxIp3ZlBBz4LOowaNujQODO1sDtXSHj8quLfYj6IJbb77yWSM2GNa9U8e8KxaqF
d2J0uBc2KNc5u9awZmNGgB9dk2rqmGSq7hke6Ac1MiJZV/UMBPtL/4Z8yzziNNpF
r8Kgtoo7cmq9oIIkLIMD/ajnlyGRyQ/sgZXLBn5XZ6bPpc9JkUsyqTLbJ8066AXh
vr+yDaN9adgU8jkXkZKdJ9QtYrKUbayPq/6vpGBf/zGm+6RxvOwHg6mICJF8SlBi
NQstSNccN/8TH8IpABChMDgSJtviajb1uQUwOoKxpmybEfGyg8KONVA//M2txkHU
QNk3ysmXbP87L1jYro3AYBqwm/SKZukFGgeolv4iu+9nAQxfp2b+Ij476OIk9vyy
c1AszTDKCbYZJ2f7y2VtiJJgOrtdo6JzUGw6DbzZwmGtdJj31eQ/pkWDPffCiuLj
9USzHdi1ircWHr/fL8mW/P1wSZ2a7SohIM+ZGNg5fscYCiPVhIUNgpTDfs0tdjfx
TVwYXbAAz0yH+lkjdmTtBiOTTAYPZWw4Nbo6KAraE7ac5ZbAZcBM7DIod84jSiMV
oJfogMEYcEiiF21rXBgpsWP6LfOmpLAmCwyHVsmGllc6R4AGuUDg5yC9QflpcysM
/NdbQiaLW9SypWN8iBrkIdeqBHDVMiVhs6PbLNvP6LTvlDx5IHhIqr0TWToYIQcW
rQi3yFm9hrLZTglD/6GqR50EP8JRNTfI+hdR8HOT9XPP54k3GW4FHyD77Uy8tJDX
uwH0PCtPJuAobFVy8ztKYIsnskU10vi4CZ0QCHYPkr9J+i0ApXSu2OzyfYps3q/T
Xfe0lY/P96XWxxjNOMnq+KEcVQO1ONoK6xe5yKmiLFHj4Q9ZIpdxgqMYqC/+3x3b
9H215Ih5EOyDwcMcHUbsCLFFYkFQhX7yDBy/5Tpw7vfzfi+UQdy54ZmnE44b+3Jm
R6nASy9jvj4mTtsZZQD8EEOrxOwGIRXPRjSqb6qbPtYkTWsZfrcnSFn2cnfEWAKL
lclDa7nKOL54OCdNCUykhHZD3V17SiHSAx4BeVvHRkQO9GW9qSNlIM7+3RoMDTnd
897pvYeTYjNDYpds/hbi5znM1w3YPcxkBV3bPSct5OB4079nnUJAPUg4hdegPXos
qdtRlFcgmB50bH9jaAu9WvZt8IAnHkuJmtaIJr4raPbUL11ADZv35XM/2Hwa6EVR
lkQZ+djT01ecqsNmfoIl+n55X2nKlRsP6Hsqcd2lHMq9rstcgQuFBLU9nl2lLfu/
qwWE6u8rK/hUvW2mkD/P/PBKTCfxBVNL2oEO1WgzVVasjkyzCA0f9aGe/zgPIyFk
5U6uqNsz/41uEVdZu8MHnI2o731TU/UfnuUDq4t0CurQbD0PBVGA3UyKSbj4ht6I
DwrKDqTB3KtGIJoyG4zUtqFxjJE3z1WcRNAHneGbmPCrM2XdoIYC4Fk/4OlrkxgN
MIZQclbW2ZEW0LNIFS4Bbf5Yaoy6nEeAwj20ev6yV+7R9vIN7XWxc8fPBkaZ6zMc
xpJTL6zNJTVwBGndRh6/e4RiZOaUin2oJEirpTq9D1Wx9tB9n8nNzlj1I+7XqayY
ROHeHjqtaoBSbzl8nDpnI256ne6l68t7Igz4ghW6QTjSukYJO/HCbYCaDWH5WFi6
fmOe8VY9j6N/3wTwr+gZsp9a5rHzny+q4141HO2ZKErTTy3k0pI4Z6NMeeCiFyty
ClzrK3ySQFs7H9ISMJ3fVflNZY7/szilg7D4cFT/asjkUv06xsPWn0esz1TYFFsS
AkKPkrwpSYFzyr2LOUbmZqnD3dH4wIhTLqFs3GbDdAvRvf3FzrV2Js6GK573Syf/
Kk+lVP02PRPD9BcjDcyS2JRj4pPnfHLNLD0mc5C4D1kHyuW4kHBcXCwE9I46jpLq
kDHnwKTqlQXfY7wlIYlBzzYVjOYRKz/UHTSPX8GMotUA/889k50MrJuHDvGo5rM+
PvkULQ/Kr1Vtmzk2XWn5CITyWAjRh4rBVUXKf6abee+jQpcMHg4ASCmaGN4uv+bM
yTPGcPBsV9HXde3hcSHG6o4MxwGkqN/wS5TKrCj51VuPFZD6MYMnilL3nqTlXe0I
75peZNPZf/Zetgg/JJAEBvCQXvbrXBpB3Qvou4Owd1AC5mI0/rUNbDo79vSH3Nja
Z1tEgGAO+FcezQx/z8xMC1/t7JGOM1Qs5ZVzjJkq7gw+GLIDPerI7+KW63qgYjoV
Y+D7eMwi5WN93vh7jIOvIfVi6GGDk3C060FTd74UsRvMZ1yv9wSGiwBseI5NKHL3
SbTCKBYlea7OxXB5coYRjx6pPoUe0bVWjD1ulO/ytd+5we5Cmh1nZHlqHH30aPgO
96WSeMv6jru5oKPeoel2IdPE2B1w3c3RCuE23v6+qrmIOmoZxkqGlq7xzVCp8kB+
rkNrXw++gSOUWAV3XzSuLq6/4kZTctCd/anYRP6Z/qJKwI/c/tqiaeYRXajQp/c1
SBMjBzPE6wm4RE21wboIBARBf95lOd6EwMkFBa59SMwDvRYxEheKIl2cXNaeoxrH
Lk86OuQQS3SzLe7+GAjZad2qhDxUnEtHyW8dYDKfx9uQy07J8PqYelSTMjIkwZ8U
eaXfS2fAaW6vniu4nBYEyBaAjsawbw4YxS875ZgLT0dkw5qEgZaGM+Tzz2odtEJE
yVcjVUkKOPPMBAP7E0mD428VaVGajiz/WV3cqzaR0eo7E9AOCuCK05bXYA3IkKfK
XvcGWnCW87wcfFRzboz3qX0c8hO6o5M5eP8wFgA08nXK3+uD4u5xWgh6rocv5Dtj
XaMscNR9k9ieSdSw2WuQbQQBec6rs6xBUR4z2YMJeEf8hvb+6xid49xrHHTb2eKC
zWEeZrXtUAURfuaQBQ5RDizYXRcDuju3OkbqDtR/feNCMj0HcYfsSWr8gAtIEmkc
bpQKQENpcy51o2RV0FvWCBQTlJ+Atd7/pvQXEziyUDBTPMwZHpl31qe8j1I+2uyf
UG80e8MtcbXobJQ+H59vPg5kfMMhycUCI26KOuNEstWNlsNbODjlG1Ex8tmYgQwI
JiYInieAwg3YuP+vBAmrwgI/WR75/zIq823LTyCA9T9W+rGF/a/Hns17R5Vj/zIa
DHUUnCpuqpM1LKDq/KzjN3Vg50ojkZfQLXn6TKBfoeZqew8kykAFtYMoIoKCKpP4
LoYriLKsD8htZijwPvuKhrqcksngX6opLjB+QWjrj3EDpbYpP925/fUWf5k8gfwj
c15nsgt75qA+tOp/zwm0s4iEl+Nd0gblbWEN2vgMbCv2DjNNljsJIksdJIwcs6Kn
1gModPuePcPx6gYji47+pdBlkUA4NL6iuywjHJuB0Esm/old+bgvWqkT82Rg0GbE
L0n/qMQYbdZJZN1905nAdNd1TCdtkIMW5DUUmQfVULIpTCJabV+3m/4hhyYiB/7Z
I2oaevcuvuXzlQWcl1GV7fYSg5X5FXy7/s9rQYaI43vqG1m/axS1ynlMqimqxZJD
GZYeopbZdc55sdOnMBWEd1/VQtQq9M1AW4dyevwTNVbW0j6aAl0geqH0raxuGDqw
EVjTLAcKuYTwhMn9pJ5Gua8M8ERk/mVNKfm6Dc65r4EvTm0s03OHJ7zqhn9iOJFK
rXsU+rbLAL8J2jFAp0Jetwhxdz+9ozdXHwYmOwwH+ErUU7eZkIX2o4z1A6ssSUOh
1svgEKJrwBy5pozLLCXr6GWdhsSPFwHso5HdNHIljtrcMoQro55lIfebwYf0J9z8
OWx/tCm/CY0AYRP4ObgHKrd+C1KljzQ3NThCcUJCneNE2UPjPXBdVSFOaVir/e7e
a8FqQ7lq0MvWDeME2SPo7h1E12pG6+8TiSBpoyOof4vqCJriOV8WaV7nwqHYapYN
bc9eRnjiE8+OMTpJQCHkfOBkT6/FN6BCFgaaxRrVbIFK3ioinRi6FswBUuX6l9sK
jZrdhjP8yzf2uIU5Y8u1FjHA4gVp28syilOMgixWoDuW94vju0Ccf35/HGzq3GM0
tZexNmtOFoTphmCtSeOOlZJyGyIesS37XhXT5l1lFaHi959wS480ixDfhm1CKmtk
/yoYNmxm7Uah6kyHp/C/AZpeW495u6/wUKg7WX2PnGJE46+RV4Qc4k2qSMW5+TbV
bEfYEPb//ww8GmI+MVuCxLCgSZBncy4ChZha/YRebxaMkPzTxYsnHQGxcXdsXLmY
oMpBdzdAdVAlk55H9N0Hgy6VGcmjA9ZqgdvmL+0u/JK/uEsIvgsQieJIwDgqTyW7
RKdi7W1BhYNnsKaLyF+ktr6rfyztJqQ8VmTnNYCQgraMyflGSUWYb4kBJghTGU/T
iGBnx1fUsQBJ6TWkXvotpNpnzjZYeVd1rHE9aDQjYFJKo+oXHZDfyioLjQzIOCGc
G5TltHXhdTSArIULIKPLz7Q17AW3LJuYdbG4IIKem2F85J/U+CslAUzFzOum0FmP
pZox2qF0Tm0CCunNPBWtAUmsG5O5N6a2mPJWIE1XBjwsTIoscuHHY4IoJPQ59bx4
npo1rh6JLQD3GQMA4BZQtwkqbOgm5cjrdrHkdX3WArB77V+zENhc67VX9aJW5N6l
eh2yGtJioOujYhC+thnRZislzHpyzyu/vxYL1yfWwnrATnCo7nfRj88jFe8r17TX
/gyp78pcgJY3yEBZN1szzhgpDlJSsLKSJ9e5yyFjo1HR+x2PHht20fFBmKUO5BRt
4pPqH75rCGLve869eu9JKnQAyE/kVbAAWnSe8tDWUJICV5kUVtr8fUaS+B366zmC
cQJcKVAMT00KdfF0cZelEwOQFXaH0ntM8v07I5dfAty4i/qCYaDdp4ArdTBJICLj
YPWM3ElE8IfQTXpQk+Ba0285pJvAACFxeku3HRURi0Z9li2UJVNx/ws5wnT+Lldr
NYvJz67VWrts63TUT1nFiiilgJqFR88I9NdKzRvnpqpTueqMx1gIbueuiFoQ7rWb
A4RvnhDkgo24xtiEpJYlFF2vkroz77fPKwN1K+nzr4qvXK814zfoZu/bLlDIVsIY
MWOwWTdOKK2AmwNIt8jqT/zTOSNYpF7PQJpIdOpSBCq7481SMp6Gu9d6Ykn2RJP0
6MOCus4bNkrWPB2xs2UPq/YIfn0PhmVls9jD4xwoPnrVGrbRm1oJ3w7ACHpJ+lK8
RhBZfaZN96ldtq1pWNKQ5lr095etxUlYx6Au93ZDAd1fznXhmEqhKlK8NKgp2M1E
/4M6R4Bfxt7ovglUqEqiEI3gmTjkCXaFoaEALo/77RFz6NfjmZmx11+ArVtcwNe7
+uQuSIEiV1dbTQ6Ajf57epDtxm0ay6eKebXXbXKjkUeeRS5uvbPoJOR0pKNNnIAt
Vo0bivLz/y/qoOnlFo5Lq0LncQrZr9bC9dLoYklmHj4sxs7UCM+YQ5hU2AVo59o4
CMBdEK0/2/vU39zXgIhJnAv4P9yq1j6G0GjDNpvBkSPyNEhwAxJUIyqc9TE80FFT
8AIlgf6Cggtk8bTnDcqT3oH/G9zrwn26lFj/qORlJdVNdj5tsKf/voROtulTNz8A
QgRRIzdXaQXG+nF2hgacNgfvr7rs2SltbiEziwCLhH97O6iixHqnSbpIKZRT+nZ6
V6+g2ElKfkliXPqH9V5y+mjPY8Yq3uAEtj1G4xG4g88mpwxfbh+uXgaYK3CJ5EdP
WShpxXwsD8GXgMaLyZ/hYFCjFpiIYEsIwnSW7ENexfX7k/YobL+oZcIVKNMAVcZt
EU9g/wyCxuBUiPS7msYpOpTyLy3j6t5t6NJpYjt/lGynXkQ9Ogg3uMmqp7XWFHDI
kdFmJRENcZzNKEOMqfaqmjkuaz6yZTYOS7OUZXa3kk0Zpr6wy9SRQ5o/EmqwEIse
FjFZPWO8gnv7jrluhjTZBdRCuApYVMFN80ZiuIg8sDckMdj1Ytgqdo4iqtKlsC14
vhbQAIbQwJnzMNXwjRtYugN1x5w5T/1cTKT/FFsjtb13elYa6vxVDUaztdTKlxg1
8r6OUpG/hLruTomJOycf+6sA9KrM/jo93fKi2UD+1nTTechAh+iUPy4+aYwmagrZ
p9aviZTZHUqxuxzr06BanuAXJtxmcucXsc/f5Px4d8FMjExk1KDMgboxCyAJc08B
2+Oe1kOBLgBhK5qhcMq5NpK6Bv7z6YpcfQEA1qvTKdY1cE5ZvPwbEm7CtGScyLYn
0lNlK6nIA0D742HcqYMIlwOrK7tbs+YVuovh8FpEPnrcIqfCaudgXP0bShOkbfcR
wSN59dCh6iy3j1ZyNahmpDT2fMI9WV5QUWL2rZ/qE3D91Ty1UToXa9qkBm4/cMxx
AFAvyw5Nvcyza865ToRs51NwS6t1dibutZoxSCd8cIqKaxyYXGxtrgp5xa4vsjAC
5+eIIgPMQ15IgrCchAxalKj1MT+zS/HQwLAEyNwmQFSzJuPBf/0o9CBkE7Au8Wx/
xdy665cxqy0dTyAhg4AatY2lfEK2ctunmXx8eAvGG7rccAlXurkFnoQ8UerecO93
vYT1ZQSK/RL6rKuI0nQYP+VUqflK8uq/4C0DNdq2GPvoHyshnZL1NtXtRIN7h1OS
lD+pcAkUIDZYkHMzBdq7SRb26EyvCM/ncm3kdk8U6laZYul4KR0YHBLuTPj6qXPs
mUvwe7sFV0hNloONQjVGnUE04j3Ybl4YnvBp4+l5PJD7WSw1npTBI8agzHkVUDlr
5eM6RH+Zk4ZzeDS9KsQX6BFAyHiND3gPgPbdBN3FflStOHo7MqbyXkeaskayfOhA
w9eozQEw5GBH3OcKTAVaGL0xMKdnexKiw1Ak5YxMCa7LBaLViFftffvpj5foTZg5
3t0o61Z7g9GbukUGouEJ56zL4N4xpoFv4vT0Z8OrDCFfQz42JtpOhrZxZIlk1egN
x8Tt5kYLBJx2c/p3x9/TShAumPW+x40Q3gx/6ZBr9MduPV3jxrlq+dcz1fActa8A
KewXWr0Wr5nGOpeQlilEyKCgdIin6WAEGjj9myNYh7wgNKV/cnU8XdgMxpD6S+lC
e2HRf9TyKtf8S7XHpB9PUMJ2U9CDAbY6ZTTcxC/tfwfrrPQNlEHUpUObXOI14Uyk
jDQl6wzmKdzGjdZchQG28VVuouqU7v5BVRtcsHyx8je/hFrjN0nHk+J3IFugIg5U
FxbIf+Kef9vOZOOEaW18AAIe++Q3vmzpp0jU9yQcfRAJ9q74tD44yFE6NNk+XjtI
lngcDsBWg2xbZLoDUrtIzcyaoS917oLSZSWFlSGfE4leoEABipBq8yasztPvLcAE
4X1GEerocTdKQ8HRGffYSXLOAhS8FeRmcLfEPfkvQPElJ61tG9ITiJpYIj5MrDd9
TRU7m/tUHfjSGO1XWE5i9DfCJad/0ID901MoQvr/mUOxkzZwKQDnTPY8j1T2FzsH
PA5E5cB7RRQC3g8oHT4jhuXte17v0yHYNdUrJubfOtHtz4CMgpVbyhwvbGEBD/No
Sxr0nDxwAU/q84zWxNS4obLQZapxVSG0zal+SlJYACdlXNlbVQuu/+1Ny2JkgBWo
B4864TzDyDV+Lpjy5q8ulhUMJoh4V8EamKeNWR7bHZiphCRbPeoSXQ6yXW59lZgO
fLOkZ3WV1or79SD7TTe7Xe4FyZnLFuawaUyse83aYthOkiY6W3O3O0Oj+HtGAEzh
zEWAxiBGFwiciEzCoYW9qfY86Pwropj83uNqlYsgli5kGERO/k7xqmB332AlHORB
2rkExHibdYPvmNCVVWWg7JzjrLlOwpAwEvNNpkb7YSgB2jxMIA8weCVQCtUHlTSW
m+4PF6oQN/HgmodMpcfmyyDapHJL9vdt23yeHWIJeO+Oi1SCsEUjzkXM9xA5mvEH
UpmSzKz1gq1xhQF4Mth3kutjP39+grrRu3hRR+CEILZAalRrBXFeduWQQSjFGOSZ
zzoshHyRjZDHSMcrdTR5dB4q9t4KeWZBGb4v8vg5Ho7BHWOIZkNpmWvwKFpUFSLh
hcFW1im5yHQzQxKBKcYE0zvv2ysx3srXUBAHeCWqo2Lpp7Uf3ejqofuOgnlUjNGG
j1j45zHaPPnyt6dDzWW4V7R7nT+Wt3JbeuxITl53jwFnnzxdhFWyEg08dABKbyos
jSUOYVvRu8ecxhk8Yo1TOzaYQoEsp+9YSPGFKaTIPOIJQCQcTQ6r6YWuyDLrFkQX
dyQjC2ZyZ+r4DCWTBg0jlSy/qk2A4pKNCYX8Omx99QOSAsZe2HirX9CAIAJcZHOX
94ycvswspZj3uyAx5EbdqKTiK1qf63jTFBpIMgfBonfwYDn2phMnVJDpzxt4Zd4C
VXjcyWJimMw5WjqjXGJnTPQ+ei189FwQXeoAhLhUGENsFgVtxxu650xtWRMrzBnt
82O5j0SU2Qnyq+7h/qkuTowMM1I1uZd6QFkR3eGDAb0Q48zzGW0Fgekyq2o5Oo/6
90RwZ6dH0U11jGSgtbgfCPgr24OIbrezJNFc5Qbd0fCZwVfjAHXxZ6Dj9/1+KRBU
m1MkXrLuwrFxY3P1RdzOAfYgyEFHM5dxVIVt+MZxtKk6YhA/yk3LdGoCC4S1SxQN
YFD+Xuab/ejIlX14fr9+tvLbVrSxuLUV23WoPbxR+u9FY8xygdO+cbULSL/8S3nk
9Tqa9WjmURnXxb7Xm+q+8evZGRSgNcsVhb07fam5oWmhTC/xvmKxv3x7bILZ6jf+
BfQAjAYh9jvV7lVP4LtmQSVTagSt0fD2Zqibb7fUL+a5eT1Pug0PcQYbd0XJJYXv
c7X0UuaC4IqNGX1+WLHD0dRDPbRcH7sCe1TAOl4KbPtXjOtCFLKYNYcNSFaDmcQy
uoJfm2cbnXjSlSAu9NVZ7+PbZnV63Fe4Qv9JGvl+5mFMLy797Uy9eOkmeuW6Nqs7
XSdTVHi2oSTS1QTlh4xagAMWhL8y/uLEU2JWyuJ61FOQwADGZ2DKHJNaxNjQKkkU
bT4OsIDSk1lp+tpCA5xvC/b7sbdNSNLK6x/+8hWgvzFW7OIABtUIiD98pV9ABHP4
7oVOxz28sbXdPpWTmZ0FIW+M3h/xPDP1FUCvq+q/zlUSdZTrWW+wHAHTRxKBQ8jw
ukd953Z3Ou14R5Dn/+SLNdMtMx0r1IciISEgKUgSFRV6TcFCgYO++Q8rTh9a8ycw
gyOsOl7V/6VRN/h+b+GY8YfggBFgU8jS1cX/9IsK92hjPZXnpdcJF//jH+PTvGV7
gAQ1/qE5TCSuHDJy3ir1zAgg7lumUclrst44LasLUW7NlVZqTRjOMpZR2Hua1s9y
ymrgpJqEe5EEHQRoJi4Ytopp9aXGAMvMD2sLG2tA7ze+tpDCJ33VFZUgA9IF3VbV
6yaSu1gqzeGdwK5O6sCNuELHmgQtH4FJr/6zBm/EMPHNUZchogUY0fAOD8lKl9/j
bUV4MtkuZYkYm815r8lLQaTaSyWFIm6tMcZfnLRH0ygrBclUbkSaOmsCEhUsbE8w
jaggehNQapiC3aZhYKlA2SMZycjHYcWzPht+alL2LKr8OX3PUnhBmWkiMoYii9r8
je5nKP3cxCONEN6QvWswTpP0WbBR0Pvfb4hxX3AmN6WlkM2tH1Id1tyeFpfxlGB7
W/7VvzGN4BKKdKn5XZXwdCUlObv1gVBZibpsyMKb97sfW5ENo5eRXACx32QRkY3B
8Rq5ZNn+TZZFUY7/xAQCjTPEui/bI2lyeudXnc0nOJ2EvmtwDEcNFmPy9/gdUnWP
tkMSf5DiDdwDPQI3qO5AHiEyHZnZlMFasv5GxcA/jTVPV03CnGbZmjf4O1ud+uY2
xiPRYe3QYb9SJPVqpd7qxEvajLSS6OJgsRUH6fqoGka0Q8Gnvl0U+apjRZKYrF/O
1mjkIu7V1eugDZzo9//2mHLWABLGlFZwi8awq2DTUNJc43zFMhVrOVObRczGnwzD
FVGp41UoI4ePX4FlCVLm/W/cZrNyea3U2XzXVLwHeL6ejY6x/haXBY/T7SgA6nZv
jABJ7rZDoa4vwS8i7sd2GZ2hpxQpNsbzQMPTKRGUWKtXkZ5QgmVMNwMs981ViiX6
hO9eXBas9q1k4dwZQHHAloS1xq2kx1Azd5rsdjLuZZiGWBobijYTDvG/A7cAB4ip
vkZOCD0un5X2+Z3qD09AREZVBZT4/ARiQT2lB/RuJJ8ccHd0m0V6zQ1TZlLwuEGM
j5KEiVyD5ul8GPCMJzGkUHVhbJnDDzzVLO2Lha/qS4VHO6rSQgPa2eXycaEwVJFZ
W30MnjusaCF/I1futf/Kc1KW8Qdy5uqGytYU87L1btQt7SRP7Up8wYSZqpXjn1ve
sn5n8/KOvpTcClmUU9zKqfNJc9seX2Hi8/5zWzcT4xLfvzlKGqqXgBXsXs3GEFXg
e9bbD/K06Tkyq+aiSs/dShAXRXsUHxjZy/ygf/aMQwqXb6hmEhmNrOVYkp6DAkXG
Ck/EKO1AS8aSxVGeINGg6Sl0ojUIhTb5DLmdPY0RbDzAmuRQZQ6HdoMV5cn+zjYT
Pd8aM+RfiRpi9OTfNeG0zhPNB6tJNSOhfO4eiBGhaN4ge+AHCd88hJ5wjVJB+3Ju
R9114KQwMgzbcflIDk6tMFGxsZrEdnHRnx0qU/nskKTkW3iHV+z/Nhbx+vuVDWjj
+ppwJcfUQchyls/s/Rl070Bt0bl+tffltV6qiA+Zdq9fYtIZFLFf0+sdyRFatd+h
CTCIQKIUOQDK4rt24kj6zF4S/8RnLoXBg5d/7PeqiiloP1p9gHMpyxTTvDZeGBfm
D+/SRlB/pDDLmBz1xCwpWZAz4nxZ7C967p5NPSVpH4Dy0fWaYLwVSx34z6nDAHcW
I+2HK0blZ30g0/THZVhj4L/sLDD6q3ZgoSGVCe2BLQUTNOwQo7Kwb8FelD9ML224
0/SZN+riYJ4L7WyFuqIr9BNHUbE2msLi3/Z2oLcS/41W48v2pmEvSywmcIFXqS8U
75l3A2o4motk2THQWI7TL5DWpvrjxj7l0OiOVe4hT7K78W87PlHUemo+pamuu53A
rhHlmZBfOSIlZF5N9Jd9jpyGrhW9s8dVyBBvBD9PxsaUC8iCLftSw6Yx08EfWyo9
/k8sggY5wgZBb4Hf419AcvuRD3B2OAa5pFfsjOqvEZ1+C79zhp5lV6yHYggW99FK
Ujp5L6bAW3m1jVAGuNkqJ97PwWuhOZk8TIyluwuGrEM/DXEpWBXUglQVHzXjDsRd
DY+xpR8Ppf5nkqyVfiChQoaC27Oq4I47nX67N79fCCiCvHSRKmRJV64OPkyknZAw
VuCNmL4Nwn3H8zz7u/3YjI8r4XAjf2H5I50UgW5I9p7ynz+rTl2Fx3RwJrreAHGw
UsV0QA5hLVb3koG99crgr2UVg8Eq8dwuTPNMjwZE+mtbhI2UFwqLiXM+M899hb+P
5Q4AQBUJX6GqCfFKK0176ZeUJAypZyOoO0D1gQiEyZB+48jwupOaZrfJ5nKVMmoI
tnu1BtyWRvuV3K0sFcP8qmrJdR88etj2LIZALTuQlifiMa1tmFQqSe2Mipp9aQG8
i56Hp89VeRB5MD/xdgfZyPFZN7eAP/RWmv8r/eqDmILZdOB2ExWdPkpd1i80j2aR
AtY8V1BMAfYNIsr5SR3TpimP5ZUmLMlUY5T8KV7gyhiH4gQ/JX0QooE9TIDTx1NB
B1YzCdAsUKDdTUUCMLW/Wh2Wnmip+J2gHWYqfFEyggcK8wuGAmhPkqIFUIn9wVZp
H3rjjoX/rHrhtBjs+hMQtc08Zy81G4xDGv65OcKj0hW496CtbeY7xgN+1z0ZYiSP
V7wNwrICyrvnhF/nMAh2Ktid3G7xO5VMuYoFHCWx2Kf8DcqMKZuHsJD4JPNPYuyg
YQZ2hrLWQLphyB1dQSSZOSiM6vW6OT2LvG8QbylLgaPYzhWRFKYF89PA8kLzF4pU
Vz00w6EC13EgC8mAzDBzXIrLnQGyfTk7TOXJew/DxIKyPG5alEuLogFlkF1de3rV
/uE1L9XTsyjh8Y83f6hvS1U3Gp7KtXSJXEgulNvIZ25RQdP2QZAK5GITE9AI9NJ+
QGMYOAp9xHTYsscYkP4ZFVTGlePgS3qJXVZ4INpC73gLsOooGtXTIFEXzgsvwN7/
oZWjGRPP8MbAK+pR9fRR98kQUOWSGX6sowPTp2lM8P1lLVm4PNaU1PMzWmNg8lzN
yO2f1QJyAW4yV8nQq+2ZzoL6FlwPDL/ODrXHAqjj5b9uVuqnTtzbVOZO+8alXgxB
ILmMFEIi0vOx4ra8+bqlFdy0dTOviVx1qLUFpjcBOK9FZilamlFEbGEjGCK443ef
q0rQrpp2SedWpTQAlw5j9/sQbf+1aqEq9mKLGgDSzjvyOVgL+L8U9biRKM9HxiPQ
OiUg3J7SfsYrWnztZr8FqUsVgbmSKTkS2SN6GI/7OkmMpmGaAUGHnvIutHVkgmC2
0NWHjd2taIzR2mRAwM9eFwb4Tb1ceyYIHcJrD3/Tyd9L8EloQXDK11/o7gveQayX
9tdc41+JEJ6feMLkdYXhJ9VjCb0TkF9+/8L3eufeg+N3D+0nmPnP2r6P5lKzLKGk
FaDTfFLA18C79g9QVtV1tllOcwl9EGKs3OU7VBmQFoMPFNmDVr/OBL2ClKayMfeJ
CjInOTTll40GFX06oV275M19Ffz3DPVMq6Lt4HPl7j0gb17XBHn4yXj6aAgHCGRF
7WNVFxQgwt7Nym+rQPgGJpdM0glke2X3FT+bU+184n6KMO9/S8IU/z0DgzgO9fnp
6lxvTC+OmT+DzSvU8Y+tdIEnSTORzddF3tHa2OdRLnwkaVN0XHJl0svJjkYQCwk3
QiCEtaknnsYS5a6Lt1GX4RND9SRcfpWRvXQLgqqKNHulkdLbC5Ar5ySdm3vD1Pjw
S1RlrOaHaeu6S7aBd0YGpo4uSxtfVXTawFaYFjHMkifDM0trR8L2DbZ5vCce9edx
tlBspBeG4xmFREshNN/FuWP1w4zzpfQVl7xovZFwvHjoYrzHN5i8VwqmzI3Am85e
gtlfUK8CBm6kky34jhz2bLEJLyZz7FqkCPA4COUiEnbtd0lymtk1P1wcUmD53gM5
S7O4bku4esHc1uZLftZPBvwS9CNut5yfEdFWw6MdE2AcYHI1wJoisRy6mEaSQ61K
dOaGKd0JRgZVTVSeKyHOD4ylfLH1cWqlD6H3mvrZ7DxbVmFrFmZLSSN/2RYoMEgg
FeZjIaGX9F1tWSMUIDtZwaZyMYAxBxBI2I430YrP3buItQwr5UWqWhYjdA5LJWKM
VOWW6GcX4Py4C44Fa3WOl4WOcCHJnauewX9FMintljLOiaJVjmzX1oXRkNYswO2D
G3akhE0dQpjO5FYyBc8LxXovDFGL5E1yXWUaLDUlPwvVJtJDPMguFYCnfvwYTM+R
0KQYzbg+zZVqINgY0ipwIsmLiejP9TaPCDwttG07wihK2wlpGMxWydYRWZOJDDNt
y4B1tyrok+IBBdlSolEWnWuxq3mEpx2M/q7zDhwn+bG/DISWv9kbXUzUL2UWooI9
QfBW+IKgrJ9dogonJCZz30/2lJYd+rdtwdUDEF5ubP0e0G+e2mkHcu167m4csFrM
gLw7GfqnaZ0d3QZT1EdS8FDarUZmv1e90qBQrhXuqmnBoVyQzM4F3rusRkMIU/fv
hrMe6f9Ny0RrCmcS8f15819Xo1SsvPB8GR8MnoVT8VlOzZ+NxlqGYFmJcpQo1sHC
929gBQkjNLV/lAz4wVc913bOQKlBrvVdRLLVcSgJYHTnDLUE6OSjrk7YeQxhhJuk
QxGZxJXNXu7vcCRMfATbgO4MGfOPt30/OFpghPjYhIEKszFdd7P0Z0sOieDsQrVm
iYoK+aO/s98Lcu+SeHh7wUJgLHVuK9BZ6bGCy6BsKtEBKU/wNn7wwDK6a0DlCc0d
0sFykybD1lmY6GZri5Z1CFPJOb074FHO/+lwRloIJkiBFdKw1Pp3DCAUkE6v300P
SrpoZXhiKczNAd0cN5dTrTUTpSVeAnpoBHoGl5yLCBLv/cGrf9Hj0027g0HTdVdM
Cvo7+rjgK63V62nBqd9oV/xA9GfTuJZqxT53zGpVpRV8zJv+/Uo/m504lopWoORI
5MsHZ9cAamt6g3akz3LHBjmMsGct36kvAiCgy6PRMuhtnvOQQ86wL3wRfKRgO91d
nnmrZp9zNH+Ge15xvbMOAjDXpSVKBVs6UFG5IAeP2bb5243+238gNeiop/B3kr5I
w9RDyqVKl0gbpXkz0AVvWC8KVYYOVyNmE5l2GefQfn59NW1oJP81Vcs09WxPdt85
H4N/GANPrpYTeOpubCrd3mqUzvM7/dZJWh/DQCUBoCuscw1WUwFd787d3Eh2Gffs
CTJWoropYwyluQ3YDVa93HP376p6NzIrw1YE1MBz2yjuEBoVC/URoMwZpa8scBL7
+BOnxbiXLjtQFdi1QEW0wrBlylkF6sstp6wZT+i84D2cBwLWkI5o1CLAR9WlIcTc
s4SPUdtkC7GSFQ3Jv/YJgMaEcwRqcyzhkGz3t63rodDyjzbAT88HhXGBfsXjb/++
3UgWUZooBV2b/lXG6hlSdrTIMY2e9pxGHdO7w16/coHmlV8ThXPT6hw8PF9m61kW
Cinn76vr/nvQbnqDWbBkDNEAaGTuylxpxCybaFpyEwDefAqorKQMs8k+1LlI21mG
s7pmfDc7X4qMAiVkvCkQHLbQLEh7hNn4vdrtXVMZ47TNlBttpWYno0roBPtRcfBi
FNWdDuLL1J2c2Ra3AcWyQefn+HtfHWGoC7jOrVKj3y7UvS9my9SxcNas8lQcTo8W
AmD0+bDdEgfK05X3fsNFMXtGHnYlWjBcEaxJldDz9aATQgtDYr4vlUjfuVKlj7Or
vTGaC0YqOX9C+dcyi6EbXvKSNmaHnkAqKCMRf/gs9T7ywZ3wBJvzNi1WPx1aJTG+
xfucLn0asCqwm9xuhi5IlqyJgW4SUF2KMn7LnEc0D5UnCkf9q1iu4TggYnISZYW6
yPh8/2Fbpufw4zMKwgs1NRpkS/wd8IGx8ybedTvJ0dTVD7ESD6DyAkObXNCtbuAE
TUx33ZjhiQB1wW4epGENst1ko/uBEQxcPWPe50nYbKMELRsdcrjVv+uasoW+O6F6
ONdaItzqHEtTAM4wB+Fr5CUGAbFra9GSymduIPvn917eKeJfjK6FdseO6vRxgu+i
OEFbB4UbW+vtxwjysD0aEd1Ge10HDKUrNVPYPsc1kMQKto4sVD1NxXuKI24wRa72
9M/xNrTb07oXpO26V3IgQgb8Csni0YdzQTdXVY04mpGmCRTszdTvb9k8fuyF5LUN
2SInGR5IHsAkPJgS2YKBfA6Bi/KuNqFcBY8HTmo9YStGfYiY2GAelKXnVRcxAodR
iLP8n1xMuMZjOyxzbut3zftgEjAxG1VFnr5Ft8OMMeKKl5CIhY/yd5ci1oOIKoc3
OgsTYikZtS5VeqXjGQLaKYZtc6wx6Z4ILUIKccwPfcLFjWzIdwd4FrA085MFZWB8
iCJvaRbcucrRpLB0bPacZ38A3DliA5DbT/hZ0EltxsxkMPWOJFYZNLk9kMTRtL9m
s1l+XaHHJ9laEPmAZfuhSxqceFGvqZ2MDJnEpeOEiftd7Vde1bpl/lr2KT5PDd8e
zLe/Z7dD0w6CM14t6wky+yWLDdrR3AWfc4gDCv1rwttA20GbzGLlJ0cdorTjb0O3
6X9bj2yetWK5NCUN19W2GMGWiLNfwHZqQotjbncL0kM4LkNtCvt0EMqnwVRbO4Kl
u2njkU4TJQcNiPq+c2FUIZQKW5JcPPAUFLmCt9cnJt62eCyjLoU+TRC1qZRlSzEU
0fYBHl0GnLtTAQDobdSjO047em32ARAc2UrR88apY3bT5sF4SxsrVTKXjsAH3IJR
q9auZCMpd2MLOLICW688QUTb6S3bruxg3DmzztK3m+JuGOUlAuDDDaHYFcULYXGW
ao+P/M+j/r4/8G1/Z9SWV8DDz+e9dn8ruRBq/iJg+/AvZ2o9hdE6w/0ospkTIaPs
UtMFfajxNEGJ/GUrEdyz+etedj2QwPOG55w5PoXUDYeNMe/lAcNIM5rNM8kBomT/
fN0qxQIeOiZ446EDGvbUpK6XTWWhc0pWM/hogXgqgJR9iCYKwYtjmVryRqpuxhQh
ZR9Ii6BbNgH8QYeKuGbt8nKOqu5mxA/3nWM0sOueh39t/iQ0gG9NhGNprUBoQuD9
CKIoPSF943GJmdh5HDazM3Ip0hxZDay2LrFLzxePDzyWOFTFQ4pKIizkbJVTp3G3
PM+Hky4W4lZ91keEKKeIwu2LbjuRoNcXiajN/nbwjevFQu2rjGd/5sjO94AkM5xn
c8DRee8jDOlLaOjuMPxXny9PimpJsQik9V9edQTSOPeZy/9PhvkwBaZ/y4Z6ShoL
0JnnUFl53lInBlsctIqPkXDdhMY3l3+rz+PKG/F84i22JCbi/yyLZPXeXLyGLItQ
H7UDXjYc9bBSzXGP72IoRCIKsyN53QI1rQaKy6uSJimDc1gsjpWvXpSpGv37s3cs
8j7dMH4GmIlf33np24sLytPBchdYR3qGt7LbA4x3SEHSBXqbjYYeLRWsCosXro18
GXb/pAHOL9raXIhn9VtStlrpdciaTcwyUk+F33Rbmwk+VXao2KdfhU0TX3flwJdn
wVjwSmis7BQUechKZV2NQ1VBeWTQ9IPfOJKiWKACPDo4izckIu+UyY88PZANLXaL
fa5fAg5NPxQgxx3kBcrGxb555vMqn/VET9Qmre5Gi++Hvad4vDQX9Zhn/zzrPATd
Fr7GPBwxUTaJ/oY3OPx03O3cizpjn1VDsMmI75P7ZBTwqxdOF8Tpj2kUl8YiEc2j
RcKA8DQcJM7Alrtbh5raK48lgyAd75V1mVlBWAlTFAn+m9372Np9+s2DJUBsIMAu
YUH7Ya336aZ3TH83eCg2Jue0yNFJ/gGtVlMMoQApiUjdvQuuSKYCJ1IXjOMokBDi
KYc36e8nCLkRvrUBE35WAQH5ttluBQOroAP5bTqg3c/wlN6isMo9DbiCvF0B0LTg
lALSiOim/MiY79r16PF67nentYNPnPa12jHGw2ChcaV+uqN7Ahj5+wc/8EcWWiMm
fo6gmMH6oMv79awhRPH4fxrLWWrAH3b9Brv69QH0IahPaHU/H5waW4eI9c9mNGGn
+XnzbNvMSyz/FD1Izm6s6oXec5uLn5XFX5aS5v1EVeuiw6H0OlWQv7Bt8Jtz0ywz
qqVG9WYF7PZPWkQTxuhbGdHap9QjZ1EczHAfe1ztubFDS6K9Lyi0pcdEdKEM48ag
zPxM2j1BaPlg6w+JjvLRXfm12y3x6vidrqk3X3KkV+kt5UNWMqnQVcNYHv3xYCAt
qD+AXPVL5/MSLJhWP59XAG2L8OYGwjvAPgWC3GpQVtDGuOTLbeL7HxCyFOo4VyPt
UYlLeHjSDMYK8iTcLmwHCa05gxVobeiZGDvoqtGNc5daKOmRXwljSmJIPjQxipkx
Kt9Y/FvfOE+TR37lb0PPwctMIebFQ72wrI18Bol04DxsH8qQoWC2pnfsDznCC4eM
xoHjGJu2A2zbQExgD9ghr9LCw0rmqpM5hLPEp621z5mflDCjgy5KFJEzUqPkvL22
KI6wRAo9h4I1/eulYidZZxpeodPRllemigdKbaWbji+wyKD9Z6tag9Wg95BfWoiH
hzRPlci/nyEnz30Oy68mIoZALBt7bojQJs4z0psNO6wsicjwfIPyqQdQ156cvIzh
0xouAdhCKXbGF2FuuxBQIyVC1S1/ZbeG4ekiMa0jRBpIwjH0VpNQEG9nue6FyKCe
D0BDUnplyJNqyTQrY7tnoAgeLfL2vl+VPLkmj1dC251CidrIYFYiecWJ3BVPRweA
sN6Bnw53wcexVJm1045LXx4oEZWdVrcMg1Po6SEI/AW+2uwE4awEDhtOwGt4Wnim
EgXeSPldu0N/Ppn0764zVLgMO69yFaoHCiD8X6NTm0aiZv2ifFKYOF4kHWgognqM
3eDWJKbCEwczUE/nwH8pTOmHrTaHreSy9WwkOyI2sDQwwvKUOSUELzQ4+MrUp2As
J2AalOcc8NulJIP8tFtxWTmo05SSiFQT9hguV9yVRWmkeQmon2EGJNHW2SXeEESc
6OVP49ahij4vB8QIV+cxQ0UCaDzX62xjDykNtbkkkbZFo2cy3Ilnt3nPkB9Hqo4A
VHhVf2gmbQzPQu5FosPkwxBXyyhZYEALk6h6zxKrJ0CS/myjrgsGJF63BDi6n4S6
nDrGyjLDDXB3nLuDI3nk/5GKUXg3Sn1ZLkX9WxPd7KuvrEDWwRfZnMltRvkPGH91
1JJYniyQs1yvVpLEInDzXqtthaRB+7ytsLa3k+HJLduXr8G2/7GPz5BTgS2tcSpQ
rj5jvH9ISsmbtXkSSdwiJurR+R962YmxxB6GscJLFBgoff1cmlpqp3YeuAx7jnJo
LMxeO+j/CPaEqNh8HwjfpRIEZXnmuf1SxiBAOD2klt8vVkJZJqo0Xkc2CsDlqpDv
irohc6u7yzSq0yHAijR39WdP7rD/FXs4YJ+vsTEsDVPvIu8AVOb2+loqPdHJPbmN
fNVeqsh/4Sj/dHVfzpADRHW/bfR1ysFe4o2qzKJjd2nVLBHgEn4RofWrfF3oGFDn
H+w/223/gY1wR9p1onjmjjR5FqprYQ5FRcAYNsciDO0+pkiKJV6sTJku/q5c2y3p
1eE/eKCVfczR4A7lAOT1RfdhOWcmbKq++CQ8n7IXV/4omfPLdPxZJGkXPKLQyetN
CYzJNLZ8NgH5UmoeL6DGuVk10wauZ8wSEvqnt6MocblFGCiL6jw79WosTY17FXzP
/xjVkBN7BwJNXW4eYTzMnQzezMpQN2mfXLeh2AxD1dwzwKTXB9dqiFZJ9HQdseT3
IaBMm9AVoju0tWqyH42MZSahTivpgGAZ07qjItYe4RZzcPXtxSfcBN1tJLxfGnYy
n9VArEZHmqsCqz5VTtwhr/oP9QQG1E7odJFACASyq/aI1GpKz6JbPYxB/1vzfrxV
kb5ULG6+eIB/W+7QZBtj8YS0L0e+sEwd2Kx/VvyGL3YXc+QR/P0Vt/u75GVf0/SI
oxC1NOTijT21Qbwcxlv4Idv/6+rYTipMA1G+ulMUAJtw5RwuDAsmGO+zxuzE0lHm
9ioB5B1OlgP7+yt/m56WejtmUMQVShXQxCzxsf2pXRU2gY8cvTLUvY3XckRbm6Oe
650XUgcO72ua9ubydLmClpeqo6/WkjEr1i8RLdKyxs0S8vXNsg7pSiUv+Ij1ozJJ
jjh6eiSs8yz/CegzCxunZQ0oyYY22mkbzNiiGlU//wJSXehZApjHK+e/1nf0BTM5
874CMz4mTmTkHPuvng2p5fCcauX+uM08h7L5mQhcYRXCt2ok7I6XIe27pRTZZF1h
zARLa3Hgwo9wx11EKfcsGFQkAYIj7Ye91uSQ6vKZU7p5iO69e85uCHsBrRv/SeKW
RX6LnUYu2wOE2RpEFUFFuR/K5lMEaXA0DnduNTmZ30omGdkQR+gKdVIED5xO17AR
4VLjks8+Ee45MFLo4K9EUin1khecvNwZmQe+9dFYG0sLjsqwOHjcbG63fyqlsTzk
L7/+oIitkM4WJ6fj9uh4Lp7objcD/1e19UPIMlcNXMr82KYmw6hNn6gD9pT6TH9m
ZzHezyIj/Gl4yBPD+Dga0oFUYMWk8vmXtKOJDMfiwF0to82A5jS4IUb67Bo4VS1p
lzr4SfcBoTLwPE47Fb1IK3n9bIFU6DHsD2IrBuCGnYTIsCqdPm3HYVilRazG/28m
lg06LRrRm8RsMk3uupnIcR8rDg0r7xmz9B+0HfsyMhZdi7ucvunJ/vEuyK41MpDI
NV4VB5HHg3IfGwa8xU0IsynOHEc706fVrFL0SGu2u9UnbOf9W+o/KsC8b2K1rlMn
n/VonDM8r3iHcWynNlS7XD5hY/hrQUyvb96JQICpXjdXn+MT48osd6DNoElMTYFa
sf6rNGdPQv9y+pbCqVJOwVEVHPhA/b889ntbVUSStbsY/6oSQpdGazcWZqtTeLuz
y2/YSHkwQUFZUkV1P1nxXFS+bOERywpBVXXAYyVU2ERItglp95VFtW+/vpeMG2If
x7yrmJ3nJu7mQzE+6CS/qomYwDznE3jRZyR7n1fh7OviNyaKQaQJpEV/WLnQdFcR
6xbxINIeewggcRhSU1HwCtGZfcWa6BKRN8cLxkdWuSRBnDEljqd14D3djiFBdIHf
n1SsoBQmdt2PiIbClR4K0yS2knEAlCM7TZOq1W07xdMDJ1+vIzw9aM/V1YcQZaJi
lBF3y6sZ9kdQ/CjuEcM7bVA+QA1M8Ax172ydegMiqptDusM1jGtp24AOXbpKLheO
eZmniyZRWpf4lNdrlHPZXoQSUa1GCV0eKrnOCyZADja/uFjocdW1LbJ/3R9S1NLK
sjdiMF631ukGPf/z2GTCQurwXLUPoa43ARmC6YgzBPrK0ogvWJ0cOlmd84izwtXj
jPeZFs3cVBXocsfkygLJN9Bv6hvA3N9K7nq+UbTodMY5FBN8b3pniugjzLYwUvIi
2BV3zez1JFKh+6mPSjl/pMj6MbYxLoZy+P1+EpuvWo5M3OvICoCdpJdufjRYHovO
FcT5EBnJ/IOLR5NtvQxqPBnCCdYBjO9U5rRNkbILQTj628LJ+BQtlNSEwQxPcTTh
JvYhjDruc+cK7f7Psy9MxG3ckKSuVoOvaQDg+OUWqehncrLxN2+WtpS7DnQGl+/P
sBj1CamJIBg5DEiIcKuUY/ArYHnfrRI1bTcAAW/xiVml5F1XEES5Jsb9CpBxqVsv
n7D//X3z5hw8HSXyytr08owyvcwdwjst+V20aLd35AYLXe94I9nbox4KMQ9KpASu
41Ks3qg1WU0mmO1jmSsQZbN+NscEaEL7Tc5N4O9KHE3ccZfXWOKgxGdlzM0SDQbF
D/DPe7Iky2z/et67Y7O9BLHKzvmRYVagSxdggHnQPHCFgk0UBPOYqmz3oG6LuSsG
2XGD2ZW0DM/blqweOGixfpl6oOCCr+FZ1PRZiLS/LnlrHCQd5uVoZaZeK2vDrY1R
gXe5i5AzanzMImbga0bYvm4S7iufO5/d+kVXZV1DBD82w2DM7keFyTOto9wMz1eD
wj8BUdYjliMomTEu9RRIJ0xor7qtICPPWa5u6swJf/UuIqL+K0oV2PB7SBO5gO+7
nM2Cvf378duq3+9BcXmneNzOka3lmFAPvHoNxfVRUzM/Fwo6g4ZDt67itcDO8IF7
0+3GUmPPE+r/2hOjWZSYXeSPHwSP4oL8hab7rNccbohX6ErRwZd8VkrCQ++yYzHx
gY8MFjsbn/KtwEpKz6veH89X79Bl6GUORqB5D2tHgBuxjGkFjj1wKQ6j8iC90mtP
trYu6q2TNd28ZNFtVrPSdNLAGtlt8Ds6nQ6EacRO7vnLgpJ9E7CKs3VTpQKoYuUD
E6Q/1bzP6DRxU+VHiDHNruiOav/sezKKhb6jM83al8EO4+yjdDfoQs3Xl8OG1WxM
blXIcD28G1QyR2VoWcTGcHMteAPbaYbyLstmM2MpH9yKR5CyuVzjQ2mDxCSozSrf
aDTrF9Nq5b5jCI9XxI/AUJCmCh0QwRgQBt4usCGZnoCoiH1dVp2vqOekS4IH+EjC
YTezG7O6wgzNR3fgWlees62zBDorUP/2XpI0fKqew/m7XWRLWRfNeJcHfzVbmAW5
iHCvjinXmnv7m0ub2fGSJrRUw7MFXmXwtVSS1dNtvteDDS4O4EjOF4QMG64fouSg
Zc0OV67UzK/E/vtSSfB7zDeaAKzkZzPGyDa5VguX9kVfLAHV8vS3+eFvHW4CeVpr
ENStGdtVtmXd+8JHvN2MhOI6tc+eAsTXOLKyuKIcKsREJCdPshFW0K5dELBkMu0f
B4SsAjllhDEFeAZctKShBfvKQFpCTgUURgYk3YQ2L+NKVLjnHsdsx99r+qnZrkCi
PHmLhgCGJB79oVaOl8KGnMGfFmo91eyO/vpdyMU/8L1Fse33+mHi3UY+qlS/TD7a
yNWDwk6aTN2DcNwdWZKq1bGc8fA5RnEVBbWS4atuFlBSQeQBfEUC0FeKcXShDje3
dhV2ZeVSIEc6RpVUsidLr4yIYCFpIclMnWceRwZRiSqH5xosVBPh++e8OXE+0s69
pBZyJSzmKa6YYXQpnjkzNSa47NuCKo3PEcwq28+dldpLF+LT2jNbYpIMcFRNEIoF
pS2hvelVK5/AUiY65u/08m2WZsHS5rovK1tyDEhrubHjq+DTYTOqSqyT1UIi2fpc
/4zVml29BgjxwSc5b2Tbzb4KXatDO0q8jXYFriUQwosXfjOOWTpeqaxmq2vb2Pr9
WjvbxHrJduGjsjXyRVzCbm5Qeux9bxYqDhxmAWshdKEVnle1w6L35M948N9N/Pfa
FHexH/wGYTBG+LrwY1/LvWv+gQkXhlpygoG9fTbk/FFi5YGnb1QH2uk7gsv4Xg7n
16CCirZ5x6XQn68DVXAl8XIKP00a9QT2f8i9wv9O8tS67lJQTuNCzuvggLoeTAAB
aKXzEuNtrx4oedC+juNeSrutq6uaao9GDjMRlFajyG9fpYp5TG+IPQTiJN/88jns
9kSVrCi56uDDnFBd3+342w2PDTBhAxM2dxIadpIBkcweQeI8oXneG10HaYdeeiO9
TY3PZulO0pyJrIZ3X4gkf2nv/xU8VZENuJ6VCUfu5hu1WOV6ktcRbr5ok4IkBgyt
jlJp935jzs3vRCmuz+SQTgtYNDX1aEOtmaHl4CxjI9/Mbf2A3bySxiEjn2Tdo5Cc
TfFFNRemI1nc+8Bmz0g9NcmS6DGkIgm6ewDtnDtKKGcxpGisLdcWpI1OsHc7ADnJ
WiowvPc1CsHIaO2moSsPdFOtSGlOYazzioUd9pfl5kQSCMkIjZVyxvQhSA7atneA
88ssDY+nbauZGWQoqSPelunM9akm+kWEXS7lUGLiH90UryyqK/LmgwAmHhrWxUrk
4CNIK/UHUznJ91qSXP57y3WjCWlVMt/Ry5WMykLgV+IvGVJv5zTy1cl1m9zWMG3O
J6sQHveuStGeBSJqF4/P1uQXvDLRJw9UT0FDvIubjEoD8aYJvTYImXGT3ZX+xh5S
iMnpTQGI5erthsrRi32nkXhRrzMuqghgVZr+AXwKV3MeysLQRwOr2C/fssobjJhu
bUzvoriaLJONW5I9ua/CgsvQKG7P89BozJjVPRE5jUVdG1hgDkY1lhIoU9FEYrpV
svzCsx0m3fJ/c3ziNw766tk6LtAqZpFSvxBUe142Bb3EGvuk8/SWdQrrCYjjSjjA
sDGDqr9zjbmmzypQv8moKnh7O2vJ9wkuEKe3M+URvnPWw9LWYIR6e+XpZrJEFOBa
Qxxsa9HgZTMVItI1RUPuyGcVFK6Ly85tyB4imWWHyA0Hp5PPhcjFuZ/y12nxPEke
kBB/SkRjfxAdecNf7A8L9morkSDzcs5VxXhfTU0+dU8HrgznGesNKjDFTdQiW3bO
0eSVTN8YGw9M0a8i2tNUYL8hoteB+DmHaVEP2PIA/JLtjTNozBQJfJbQVwUksbKz
l3k3uaxsoMysa7CR1mLQkEojQZWHJaOLvsM/+wegT5ShzWhAYk09yDsV+yEDowOq
puGG/9IbATigNYlY3wqxI5T3aIe/XKEwKwuH4ApJ+wOGBzceRzirVAnSGqMmMVT2
Qthajc5Ot7W3S/sIpGryiW4aPSMRv+kfNKHBTDQepRDrtw7NlyVzDgZjvIZCvbeD
4BRoEscXBRfhz4/Ev+UULvZFuyCW3mpPLAlZGtPqIBuIN/NolOu5YYlgEvaEC+OF
e8+kvD56XGtj0XYM/CjhliLDvquVdbyW8ef/iH8saNUxptfgQB6S3DF+Vf2B61tM
xRcYdR2Nj9GjyznfQR3Wg7i46nRkpcVeFDZudajwFsH8cXtGtC10or+bYsRJsDjn
KONJ1ouJRkEJsuaDnECPSWmKLGeHDKAejWXEiK5SS0NgDhUqx8S1IPEksUEO+KR0
pxhkQ9kH7mvC7Wo6rEUQHFns3UDCZQkj1iP8y+gUoBu9CeQY+MddQXZx9WfPyxmU
OdK00ifJjVvAbwrtxmmwP6/+NGNGcjKv+bXEgHMmQ4/QZ77rfvPWgL4Z9vpesLot
OOYQeS0WTQZUJqdE1016R+vKHjo3FDtEefifsTklDC5+vfrOuU8h4ShP/SZxFjo1
18Ev6sFmsBnAzIHfXEm2njhutwAq/9JU7n+XMpFAeRr+AHLKxHQqhyLmavafv7FK
gMJremhWFarT8QpB0t1uBdQPgSYD8RwwSBeELZpv5gYh/dWXIn3ylRJCHGZvx9rW
njqROBZvgEuObBEetQHJJH+n1DE25bfznAUX3h55FGVhKAXiOlnRgRIrka01yhBs
Up1H5XhkDxCepJBaibCZkSKTd2yJi3GbMhdNyw4XGzu6Pig/NhNjKKJ035dBnFaQ
4AymAy62XJlSneSo8K2m9FfrJZDFa45/+ICHqXIuQiEbaUDRPtGD1/Fc+7z3qYaW
UOETnFVKHR9gTVILUcHi31QavRhfUTiRGcfjTNZRO0hW9DTxFm6hgv4oJ7D7WkTG
+ZiBP36zQhRrQnyaa1MDv5FkPfjEdbgyDwExdHCD0WyH3R2G1nRScYWqowyLY16w
NByyBVpomyHWs/jy7ZwssnUvS6ReYyLRwrRpLcBtVJhXCpMdIa/Ba7/rMdlJlC3S
2MbdeqeHcFxGU9sG8umt3ljRmH7orWtZfHH52M1gJkjrdT38/RH8ZS5asC0u78rJ
a2o3F+YG9/+8JzvTVjNvQhPqwP6Qei7t567D51r5NGu+lobmd8c7Gr2GvFNy1luW
ybQ+Ptgid7Q7tL3gXy5w/jTLPfFxBnRxM0YZNhtz/1CtFaDc2jH8bENol0VkaqRz
kKgNRG+lNlFJQ+q/XIRmd/LO7kW+k8Qn8UDv0TxoIPLBeVqvAT0UyL5qbyK7/6Yn
kWPLDqc3vGy8/q0qryR507IA7RnsTkseZvZGG1hFx7Js7uZGAANKZXD0wTqYMPTf
Fz6Vq6Za9xNqe8QOVAYXTtKXrLec0NFqnoCO2g2Zu+sGqLya5y6Ll+U/1fPU6rjA
llnsL5R5GPyLAHd/3HKx73Z7KuXv9kBaTmhJS1bmZ7bXjU/wTLwZWKHl8/WN6fXL
NtfZrqdYAUDmhzBrU7f5LtyAbowg0b9unb+89L41s6CL3+qF+1U8wC24lMtBL+kL
4zTkKz+vB2r9k3peRyIs8UbON8CF1vepTwuHRuhpz5phXptHkXxpNjclM1gH3D3W
xuDjJLwcEE9PLWVMGoTHat406VMzbl7sVmBW9iM47EyTEKyDYv5nEsRQdfMt8/yj
8BzRMYdPXscl53fKv+fr3HI4oSoCNlPb3faWaKvzMsIRa5UKFzz6vdPJ0i6sxjh/
qcXuL+bxoKivt7A/srrNc4kCp1zpEpDNwSXAkYvOb4OxkqyD7DJ7/bYodUB3A1wr
Ifwt0cR3ZTgOMwbuEcr6YQ8ccZKh/j7dxA3/NEfl22vdfPh4Cauyc02F6UrkYOZP
N+4vb7+6wrov5dEWwdwQVnI1qkyv3dhRsqSGV67QzgcITqG++LwcJCHsYxa0yzAl
x7q/qrVGAVJfpsG8Tv0l+xWSuCscWW+TuGuTGKZJ0PLrAR3rri628krKJIK5cXrN
LBCRoyJVnjCuxNC7G0oii2dBpGHphV7Zd45qgWde3Gn2JVLm8hzWAkate2WunwzH
qW8kcg5QvU9Crx9E3Wlsm9AZKLSLNyu23nPEv8SxNK+hP12G/P3nrohyJqz/tC0E
Sk6TkvKNkdTW0whGteN/IQoL7LX2QI5rvSIHI567ZjM1GADm+/qcUhfTq2Lzzbso
RDc++CD8hTYo7UKMTz3m/MQpqLVzhCCVuL5mjQiedjbZtWrU6yv4XniKamQifPNr
NBKbH9G/sfDhkwY+NMYzK24xm4F5L57c7mBuQMtp0cZ+SJWsHpHDyF6XmGl4Blq7
sUI2YTR6x6QWZEkIvkFnEbGC95J7FzTQFtWoE3yikA4cvt1GLLOa7EKt0HbrCo63
m8R6faiT5szK9Y9047pAXzyJdIABRzfmem1GdVX0v2rkT6PVDB7pBZmRZplxH045
skHmQPo1E/Cs4MnfBxO1ISnztsEvvRiLUDpjLY1SZRIbuFNvJnZSIsD94En1ZY2V
kYlKU4bz01x9qIUq97+KKFITQQI6ghPYyuWwKMJ2DW+xPellRrXrMf3Z3vFfUatk
aj8OtWLQgis+wKjdSLtl8l1gjMoSm/6sp2JQlq7YYLv/xRnKaasn/obAR2aSbwxx
8CU6wsbTiPq/rnqYeLKlKNeORMcEUGXUwcMJWwdAPSK/PW8zKy99zmydfKz0wvJG
3XjLgSDmS48+iM0lmzgFIT5ICTsaVIDLMMCtenxt8AHh1dnOtXmtb87hFRN/SKGt
JsTCzhg6av0lKpnC6/jqqaR8RXsX6003Cyywk6BAOPljN4xghQwobibkvKsaqRIy
dZdVnF0urZd+LUqlGbC06/41TRl2ZuT+MRUKxXEcBULAQsOzAC2zNxcrLY0KjYk5
oifTl58gzMP84dd3xx2hLrhPTxdzWbU57nDekBh5/ZhRPQ7a17gBpd7bQF7ZJBzU
Vp2IY3kjdc+tKwb7rWwHyyz1M2lW8ldKLUPdM3iVjih9zJfr+pukiebhFAWeV891
vQfy0bhpoG7s5Utda3e8LSdiWFzzbxQMrwTlDIUrgKbJb+Z6g5OaZmAYOur3s5LT
CmnmuW6gU1WusYR4MXF/W6h4V67aUCZ/+QutrkpcdjazlS/h/lfpIZ0gmfSETr33
9JB+2YCopI1FVbiLcP5YEXmoMU5WReykvlTEeqZ3NZrUB/60HT70gf5w5+FyaWOL
oOFFQlWnax+7tbLB00cogzudwUnN5vMIFDiJ12a4eoCimld6oPWFiYebNnEXLcxT
tvKsSjfXMClSfaidNmSnBMvWm0HhpSBVmQPuPlg8jc+n70DaR/5mcgxVOYjXV0lx
0Sa1KNnRu7ZgFiW1WHobo0uqiYVQVHH8XgFrpo5SserypLMumrKyLCVLqfo8jYg/
nY7VDTZEgAkBDlG9/dGrk19wI8FOTBP04dz3FhYPrI12RXMxOjpy0JMAQ9GVdCSY
Vw45Qgkuq2Xt0q9FlgD5kpFDO/JgLZiVgzdhI/gaNpgtTEIgdyjIqyLc/4kGzbf5
jLuCob3WNDS+udOMOzQwG1u0Qi25GilNFfSW34l34SADMtCzkbTGLH+hqgqxqCP5
3XnssEHvF0LK3g0BsxYOZa7lx/T2NXdYKXz3ABtSolyiXJ64q7v6aYf79MNDS6Nw
dp+DsKHLPyh9qrTFDUDnsXBKR6RYkxBvxf6UlR2Gm+l9zB7PAyjsrP5o39ttG/M6
amkloED6sThtcZVIaUqgQUpAtGLJ1kddjOPaGYfhOuvVBL0jX8fzQ8TXhaC+fu7K
B5uMQbU1IG9NFp/lrKnWOYksd1U34MhWKupjwF5fcxpriCHX/GJXEgu1ZIIAZ/Kr
3X+nQkeazfY0DxKCrBqXYK/S5mGKfRgaqySTwGGmjTIUFH8IaSbTKzF4CQCTyGsl
soaAstA7zjALGXCqMQvV11Paf5itfSJjVd1w1QMUgZtgcYbknrUuqyAwsa6IphQX
3essdfmSKKJrJO6+lKRuZkQ2/0jhev+x5NiSu9V0V/8Bwo4DRLZ2nvzvWyV7KOvB
u6TVbe3YtBmqnXAWdrA1sT/X7Btvtl8Jql3g82d+Zlw39T8PCjfmCC07Nl/8tn0R
jZh1G0bqQM06XnGjTv36NIyaUG+QSoae0MIi4Iye8SUPtkTdwj0yPnHJCPWi4osx
4EASaLpDg6NT2Eypzyjj82U4+4hx6fR+d7mvbux4vO9OcDWQ37gLx6wrYEthTqfm
OvGvKsOnjWWoLuySqLMnDpdSpmH9iHztBrwbxqOcSi3TwNp2GH4AERG4WSANh/Nf
beu9ykkZw9Mktv3hgtY1QyzIknWO7BDbfAiCYHodel6b18xA6WJl3WM3l1RW8AR3
Q7V4GTegzgcuNaekB+V56uPh6UWSuvj0ey+d04bLx8Bj6jb4hayMnBjuLzIpAbGW
UEhRqwamXB6xCsZhzgmMieKcYI5svqeML/ecfKEWY0vgxyps8kNmutk9tKBIgXS/
tbHdQBlHJhwTAPzeK7m31V2KZxDXpqaJLdzTuSyiAJt8ucstHSwqI5BelRbJbpGP
D2WDydGYmKSlCzfyXBHSmd453ypQx8Q6INIyJZUKSk8tsTnHLKsBiYWK7kf1eSqV
0fngjhyDrugSLurVmmmYTM+L5cVs2BkQZQ8SDrDNh2Ai8JCNqgpIWRF5Vu5RvF2u
4e1GfhsX0+a7Vo70UhBcSKmGFV1e3cXwvN3K2tKmC7Toq0WWORWDKM67g24r8oon
xIaJg3KZ/NshzDO8y+oem8MPLp9+nWBnU3UhQmWFcKaunEijruzBWdxFRy4A8bR9
0XlXh6XyX1me4Nd0+B5KKUVmEsDGLCz6A2SMLPu9fqiRny1u44GDw1Ndbg+jaeGb
FyOBxa0FW9K8B6croCb5F4YFjeNqhfB9+528n36K1sgPXqEp+RYnmZq+8/+9BErs
SAyIUAjOde2rV35b0skifA1vPWDD6Nq6FTK4MJFwe3IqQpOLptQRhHEJrwFeFDa/
XUsnelmrU0gDvustzRayOCfG/9n6+urUx0e8JNXZrFB/Xqa8kpslnE8esC8s1loY
wn7jdJ9i+WrUUrwFX7tUhy4HCLSYZjy/YTOWalYhpqOQkrluZ5as8IGPS8ZtQNs8
0fcU3m+P2X8OU9sRdt5kSbkWcTs2Rcd4vgY65Gb/sZnCznmmbzeWq7Ql7YvQWiH+
V3R1GQZ/D4PgLgyfWLyiZP1leakd9kTiQSBvVEdcrPvPKmsYkQDrz9E6eiwSy1fu
eg/3UAONHk54s6z5JI3UjFuUOeOSpMsuUwtYG0IakQ5F5Zoy/UBy0H5yezVPu8yq
mUIlCuOYg61YIHCZ/Fvk4npZWBNd8lRWgKqGNyhIiIP5kxx6TbHI75Mdtq9jrSM7
ILQF4eP5K3Pho6QfD0wxQcATb9YNJe0P8T3/AtohsUZ4w8NpcSZH1lrJLB27CSiB
KxNJdkbrsTiN6ugjPyFpP6GnTkoGeyGwjPHHVZcO7AuCWbQu6kmKI9p5r2D3pcCt
PYCl+vj6b6wozuuMSJiSC3KxKrn0EtTBmGCHjqEKDDq9VeW+MZeq3lZTZpFcQSt+
CtgcWqXWYfP29khuXCVNHKXDrSjGPGZdcW4DtVKyeMeA35ZiYiXEx3wzzPEW/Dfc
nShW/U+c+9fGl8uA2lWVbuLsv9Bas0HedhT+1erVMmrX+ivHwLIsXX0VC9gu6lDf
vHIU6uk2Z0xZ+/HP/FCAdOymSTQNzvXWKkbNVsbq03NJTNnNBOO9r2y6qATX+ef1
S0GvkBLyT5KHtVfl4NRNdWKACo6EDEDbPNhDTLn45wIe51v3nBNdypYAcr6XHLBf
NxkHuKkJeqHNP1BdiL/J04CXkJeN6L1C3NmE6eG8RGf+sQONs/Pfa3aVoJFY71sk
7XUzaUiHSckAJ3c1eYadU+LAjh7Vptmb+YoPtTmCbk/+VJgXyb6bxkvb5B7WK722
NjwjCWgSAUfGwrk0YrX4X7aMFT+M8LUs+pua74NxsZRnp3jLWM1CCFD4eU0vO0W6
uVomxIcyIX4C3HvudCM2bnHGQnN8JpURiTBYuBP6fujcu7VJbNhD0CMDPbZMCdok
EnKoeme6z//SwS7iqg1pnNx30crepUBhxIA36LD63NlStkOCzFNJen8IHwqL7KiT
b5cWx1CO2s7XwjlR4YU5fArgtmcl60RYM5XMHVPnRMD6eiZEoSeZKf0uaNlJ3TKp
Cfhi9hXx/uSApCtAPD5rPFl3gGHxR/HSKrvosJx8/MxjOWbmgPMIYQY6YU1zYnIq
7JfqetT374S9qxiyXvo+N70wmYE1p+nD+XzGjDG+0xKi4eix8XND0Nt0NlpeXoHI
cUmKSvU6J9UZcU0ERcUI1X+MHPFSoUhsqtsFG+MpQOgBX54S50WZuSRzh8C221HZ
k0Ek495XaWPmHhCWcsrw6J7+1KxthoIsccHi3zx38YKw64uurGgYe4/DlF9nuyFn
vkbaEgQ/VIMpo9Bo4z5KI9BZXjL3zSPvEQ3cBXBl8GwHl2FenMu89gj5stE5uL1M
U/3Zwo/8AMsz32FcMFsKdaRiKS1fH+EifkURtvkZ8iGdU+8HcTs0QhCstM1R2WyJ
mCq8t+JBl/uk9QGCNNHHtr0qA0GVvNmhNgSqKZLwzMA7nS8K89hpdAo2nRIwRBzI
6+IkmwKIUvxHsusPjuK6LW0yqrQU3c8KHvwT1sHyZu6aR9FAp75TDhTlQjrQcAdV
L3p9KNh81JAfDUjFVe/N/B49nbonnotPCJkiFvC3mKXZvlDOPM5XvjDyDpBtGp0t
lBk7h7pdnD+62cGyJnXDUBcb7EuPmqzHG383DuIshSZEwsqjbYl5HD/fQu5ScXDX
90xNNKkrtVOwEkTurVffsGzUthc933PAVDIJucsEtaAXR511Kll2y3TLkjwM3TdO
plFeBPfFMDGc8IhoBUSDrTPs/l+geSQfvoyvcEVK3Ywdqx2DXVmNnGPK1Lq+RmW9
cHnWxx9AWPdFaBPVxePWHZPigg3AnVigPNycj+2eF/y6iUX56Wt7b3duEryRLkqW
7RWrAS7Pq5AWJiiC2AZiyJwX7BMlXqZSCLHYjolc8G0I16OuI9hzFCnt8U6Vqjk+
`protect end_protected
