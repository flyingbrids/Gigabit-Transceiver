`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
QHCxKTjsbXl8yQkHcVZCrAKppIf0IHr5WMQbMMvCZO2/kxy5nhb2duQxUC5f+sao
CPriezlzJFhbGCZRl55zX+XUgtTIcQOywW/dy8m32SdaBMy+kakDF50QAQLSwrhB
yqfwV43vdzC5YQIxUJwd2fN1DMFP7XfKbr2QczCgstlkFn5tHPb6bqvwQVVztxVH
rpZPpG16GoMkoR2tP5RRbFSJBL3NwauR0O62PPTaxO+jqO+QLWEdz3GQKcOe5u9z
QcTeLIbWlLg3YsHjyHEZ4J/dR+n7IO5Rs/D31wcZMhwgBSIqrVT4ilueOjLbX+IL
zUe6loWJSjDNrNDUJO6mMA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dZvVKnKwH9LLHKnk9UP0yOUIAEzPTS1nSQja6RJsuk7Z6m5XyGxU34euPX54Lxkd
FpN7r0M7cZdBFyqkvIC67Bos172lKH1/6L6e00K+CkssKFFbFgz8fIUa50rpdU2V
GKxDzz97GoR1ccnSkLwlUwvHQT1vwGDik4deJKQX1sc=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4064 )
`protect data_block
ko+jhBvkSqxuyoz+RPZ1ywBMUWBccyBF9ipKnxV3BrxieS5kbKWLmd2HTu5YVzD3
kNEz/NLtPDA/PLT3/zw+Yo9aGcKAPGoxjbsqHTxF1bz3sjxjwqJZjmC+kZV52YgX
WQdVNeT+Ns0Ln7Kru4Q/kkMsvZQ6KqLq3bryljG3CHmx5bnb+q2AE9Rhc5L8eXva
jg3hPEp3Em3OTkYpqh9kvit9wACNjhW7uMK4bEOgW4mB5UYZLyjEYyjdupzaMhXl
zX9RCUW/5FZP3dheooHapesIWe9JxNSwkqDxNvSbL9zjFZg6BHXUUnA5C7Lb7kBf
TWGJplZbgoXhPhYlqmHrGR8tKYP5ki2N7JWFjtNgOm0Br1ri50qmw/Sywmxs0ARf
XIlcD0gHU7CqwUusre1Yvpyeeukdlfi0jLrf5GG8UhXzL9XDpr+meuVMOiDDHXIn
Xjdv28rpMuGCWi6G0jLliY8RUknw1ZHpg3cswk9LyyXSU7aE8Si7CBHpW/Vz0qIv
MkrMOg7oxm6mpCcn+6TrhrGuSWWlZzE2AjrEh+9u23y8RVWFAL33+PX/CmOAt/os
He4dzgKxwijg8FtW2AqhtFyNH8IoZRtl8NfRhU07rLxb759zobV7rgy3dVO+cSkk
2smpD0JTX4DE0Q4TjCUDihIaief28ldZ7Q+gUFa9GoAfvZylenrtJgGfimpOOLOI
CLpKaRTBecgz291N9Dl4Io08NIWlW6dLvyiZgeMOczMJCD3rPIpXVPQ8PmlBiVDz
IXWhtdvvSZ1Od3LZfgz9Ni/B+B4IIulJ2pSgNoWnRke7d5skMTnPRSOruDISHiTQ
kcouqBDNMHKMZVcRRFZo/bNgo0uS9+xsAgVrVYASKl0s36zCYoW2tZklCuGq7fDU
sR3das0FRMDutbfUsoGPq3COavECtzxbLoO0QDNas1rbW3I6if9BFHCQd2zlz7g4
WpTTpifGaDF7av6Z0MOPq+ENzrZN9PL0CA4bHFnqz457uKE4pnw+CmJGf7Yz3+pq
mGGLVGSWaztWUqDkb6BYRV7R84sX3acF1Sd4A5f818JWEWc/tWzQKSuBl+tHhubQ
9Z0CLcnHj503FAX4iOQnvHXR0dEtcm1XQkUfTJq3UKfyP7d4pKh7jM3J0El+lOZV
WBXqOMjizvMROnQti2zRjzO3jNH8yNOmNAeV0VI/QuHqR3WLfiIhw0F/yOWeHNI+
dabvFvrA4xHTSbHhXKa9TP2GUdDD/TWkkZ6YIifchdyLeVNxbxJkJ9J7uvhwZZtE
pggqq2BLIsmyD3yML4pMQESa52+WwY5tMeQzRCR3DcsJ1Cdc1mGmMziABxb8QjZF
dWVJz9DKamx0Ha1CK962We57uLJxrVrXQG2iFG3E+QwFPN7aw3aU019B7+8HxX8x
WruZ2lbZEpqoWFeUA4PAtwVLLjqpN0LGyqw9gacJ5VSIvaGp3TsOlWXKriye7QKi
TsG7FPQQsdQZkJeVo9az+X2l98oCR9X1gTFWxE3MgJ24bqm4pzvOPAUWKOxVyd+J
9EEhbXr27E1dGgnmkU/tgJVkbEO9HQ4tU/dTz3HBWzzKA2xbdEyx6/C6/HL6OdxB
MjKEIWVOa3DSMVm/kifHm4zFq6b6uzBt9ns3UWqNLTMgHu1EsJbEpeDjKBNuzrI+
UxMY1PZ7W+uoQ3Ny4BEPxJe0Y4Oo9EjY+sQl/qithm1gsRtqpGddhYXsgjAiDYIh
sPxYzsOuh6Xso7jwirK6JfkPzpgrVG7YcxTemuINu/5Gu5VMar7hkZW7VBf/1fWW
qAcsYvL2ewXEioELbqeaq22nUH8oKAdOAzpAHMQZdZUnkVuCjt/7e/ABd5gL1ahT
hQMFd85X2uv4OC/hnMM6dQONvaOWWKYr53X/DLgvwmtfWatqqRMhGO5K4+NZRK9q
rJXq2fapaV5wUqygjwaQ793QIdI8RDPLcRkwPePFsn/PUdDOTmh5SWRLUlWzlOyw
WisJNEXmVRclB3WDpFJi12AEsekYpEg6vze6IdZ0mOcikBxewwvUUoOsDxvOit8K
yLOlp1f4uzO1qxdpoT/FJ0RiwsKrSsROKWIuHSj8nbBOavFZwSdS7MQp3iFBiDxE
OS7O0Y09oNvss6llG4VKtZUXceZrAoRVlqYPYsKOHMc+8oqy3x5+4v4mH8J/ZI4R
KMXogmRc1BHptCw5rIYG9N4sHhx97zOGTQUzBZIjRM64asbJSxbCtfQeFsCc8kyj
IoOLsj+HtWJ5dGktiw3w94E/HKk+Yjf+CoLLbIJ+OhYQI1HJbaFbUf/aoZmSSu39
LoyDKYCjmCOZzY3oJFFjxA1HhiB+wzrWqHGcH7c34v50uJY3Ipeha209SQy4CjvQ
ijGHu5bdtrsMZAUksO3gvz8lZ/uKxMSTonjTijA/B9huWH01ui3zD4wA+YNT1eWy
9KyfrA27CPIXpaGaKA7RvA6p72nNDLi+l3zwIMWw8VwiDXxDp0fjSoiBS4DcNNSZ
u9Nc4etDVf6uvgOxqEsM8kFW62yw9Oa8P4kgXAd7/2dRTWivXEFogAG0BpREp5kN
Nh2wusWOlz2+mqgtFnlqCtgfplT7HXIYWE8RKd6J1i6e9D+DD0mRMC/XfYUD35xJ
dTWVIC6X9UL6AlF9+n81iHyVPOzWTe8I89G5fura7swHEkZjdASH9ttRcQ2nQVtd
2nvPeZv9ZK//RtFJiKWpzzhMx0c+0G9Kl40lLJBmxh1VYnLweXqfCFp3/ta3PEIG
2rbAyUExEb6aqQnHNytOYDoaVodUOW1kKF624r7yP35i+6mcHnxZC/rMn3qMZQKs
oPKPIuI7Bh4kP0PlAQ7Yy7WtljSNEddlqD6c/blByNewoRBQj+GvUQHx8mFDZW8o
4gMBRq97uLjP9Cbb5ynu5I+D90bJqlutvysjy1hVn4ioI9nUiISfJGqceXYtCjMN
P/vxaIFqwaYhGBYJflNds6aoqeTasU6KxtXjcXhHGn1DJGChXjyycV3KKFNcABub
fDuq9jU9yOxTAv+gPlOxoyteDQvDherdZ38vZLM8njBoK3lzSeeuJQOId/xMgVZ+
7KvtbMH53T8Tn/BuLtMxLsBkzNMtcLjQiF1wqZqmOW+JOHFiR41RtPBebpu6WCKy
ODKzkrPJ6YD9h6Gzp2tgkRNxph+OKS/tww9rQTTN2kbGLkmpcak4dSOWrvhbRa7q
HyOyU05Xuc/45vDr9hnVDQB1/Lrb/ytBJy4qQnD0vtdgfLEtF3y12VuasqmOuZgQ
iHYzHkwydSrQY7bmG5smkDnQtlaqVdGxIdI5ewx5jrGwAuWSlWBbFg7Beuea8uLn
HYZo8ihmtHEOBmz5ijiNHcDKm+FsdaVTia8YFikFOtjk4joOUrzajrXh6s7fCo41
422KZ21xL/HcGJ8eB8UhBkPWDykvfVBkymyGtKO1adV/GO1EWRRXv11StsPZ6+MO
iMofVSppayBTHVrMPVBwBEB/Bbkk03WZU4URE8XXEpIzD+xjMpB6eiUEINp62UcP
xTMaEGgfGCEwykNMwdWpMAk25AbApZ7p3ydUaZUCCGZag+/OPlY1d/uq1I1a9ZnO
c+yToBcJ5L80hx2X5ejjLIAg7XF/7oLepgThY5f/yPb+dgV/uPqiefcm6EjV/OyR
2Bsawy5DMjHdAEU3YvxGxAtxdFsPH27ZQNYjeVZpKZRRBXRzDE/0bY25cDg1MwxS
10BZXloK+a1FMlpFbKcdWqKqXmV6j4IWRuR5nn3BeEzuyy+4FTo5oxEglJr9zI9Z
LToc8ekcsHM8d63+i8S+KkHsbXyLWQHwDZ7oPqNc0GtMhXaw5GRlBg/oWPaBAbvC
a5wAYLuUBHhQAzO75F4NWRgeGcnNVSlbL0vaiXzbaUxFmOcO8QdUJdeiOm0oWDaJ
l1lDVGMcZr/BBJOaQcR4C5uzyFYck0W0AXnwd6arDjYCP6o5OKdgSBMZ3s/9O+D1
Tw0hE31+fwrPJnpeQ9Ql8wumjrALRUMbbq1gTjRcJ8oLY6lvET9jkyL2aWSGRFgE
lRtgVsfwskM/YyoeiCvLQJQBjy9fHEgRkVdWNdOLrW46pO3ymjgFxEUbFCJ010vZ
GEs4HN6q7a6CiBxnH16FmMZRpZQ8snk+DwtbW5VkUNLJ3TfBXIrXuTy2AH6fYA1j
sGi8MWD8BQN7RxtTY31cZO3JBQxkyLgj/vM8mdL3UrU1bkiE2mwrFCux42VgGQW4
S5SIvWFAwR1g/S+NJ3fCDrX5EPlTDyFsZj7SIZhLEw8MJBZo9dakUbioz60/C1n5
A4Y2eGEghr5D9xrTocPVsN+MjEE8xNJEErMojeLU5zFkxfqEf9GDtu6bNx/tBvFE
z9BIcLnd32MJ+LJnV1zOVyhKoqnpgJ0VKJn9qlKIXNSl/VudUl9BC4eF33vvryAr
zDTT2bxMPKt6WlUtIZe99SHzOdfXZdOt3CWufFiD8S8CJ24VsQ6ZCr0slOAEZa5R
g72M91TsisvFo1nd8QEC8CklKAAXxBY//u+4ywIdVpNltpCdDzvdreR7446keXPy
slCaHL3dTYUVJY6hTUwOC7Uthma6p9iVwOlSwWtpbZSI3MoHOwWHpIaUJNJz1nbt
P+gpvTR888rb5ay0i3YrxAhXgS8u+fq9HqfTWhRZgtqWuzXrnZ2lUTPBmqvXS3r8
X9UiXahaMmGc0wXNMS4L3C5+lzwg45TXiQm9YBMYsR9XidEikp8ORdFzg7qvX3Yf
Cmup+L5hMUCmfR/hIBOacQuwvLQqITL+/xU/CNXsYQeP7jHLHJolaZUbTyAUj33N
x+7G8PqnTU92DH9+JrdZOrUYRHvUcI6JQPgkHd/I/6nUa62+ZJG8InMXgC9OUw/H
6hP29gIMVNKzvrmPDbXxroKUFCKYPDiiILrHD8YIjJ3yUT6dTHy6dGuqrxARCb8p
tc2EOs+apCrFy2KHKWJto9+Lgdp12kGXeVaiBmNtfIYLF+BYJDZ0hUuPyhawg93C
sAqHUuotBleU8gCX7ENvdO2xULoRXD6D1WirxuxP/VfWL2wSaUR5aJ7uqYZKmCx9
D3f03sLTDdUzGOkAyc5e2tiUJ+Ehyi/tos6UXpzB7iGNSPv8Wm7SMvlLCRm7HMMA
v7QMrEOtX9mF8N0pooAb5fTkrOsQAr3oWYqeX8p0c5QBUAk3RzJ8K10qZqugW3Kl
Hwdos/csKJLSVOHbOZ6wPawJheyYoVPjF0+WFGquiV61NbvTS6dUo694leBIA2JY
p+RiMVCUZFo1hGbrTZv4z0KmeFppLNMO/YGvBhEDtJ5v+JY9DzFWD+ufWZutVd1O
nOGlM7DxNDdynZLgPWtJyOqA2WFK6dKOwG5nmmg7IMrql4rLO3tuGrFF45tgq3T0
RKvzZjQp5UbewGgO2mdpOMGBC17PbCgR5VKp/voOaJo=
`protect end_protected
