`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
R9uZ3J1qDKB2x82tmYugZ9kyUcSo9q4oR+WOQhcEPy7JIJHK/wX7w+eoCLKCEQ3+
S+lGbAbHibLbp5BTNkXFccrWKDcpOjr+u1+l6+TQgRuGrvyfCz6+V9Devj86Cm78
lsBAVuFwnKooNF7vbiIkrxx7HMQGpVxtRaut820TadtR7IbVbl8ixz0+T7FOlJ4t
935PUjFe93Q1S+1ii2dK8kENkYVD3FgpIOX4Qhop30BIbNoI6w4aLsp3A2zKmt5d
iwUFE2daFID8ZFIPKdEKmo8kOzGKf03wzBxKVbhsHkZQjXxQ92xVxU91cIfVj9Fj
9+fHhze2lwFUyx24B0Hnmg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
L6CNsgzLGJzBu6wwfrqqwWlAEPoAR6rOhL3LPcn6/vmAc6my4Z4+QVL6hmBYJQcg
g0E4Z078AoTJe1O+KUWMKzSw7BIRnMW48dJh5rjsAnnDCk/vgYVHKus/bRs4xvCL
X9RJouCwwj8QsScGs4bj82Rl4BlJaiz+kdk1H6PuLfI=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3664 )
`protect data_block
dB/YCsFpOAxLXAXG0P9WuWj6n647+COnH1FQiZ3OcP+js4zppuI8Ay5sISPUItcH
hkRCK9q4zSvVVkqiIEpKgUEOEfDbxx01rQ7OY1Ugw0ztT65JEuDpZOx1An3uDNND
32bmoiFajyO7gLOxWGDBp2WCS3yEiiBPG/yfXPiUYtVLm6EvMu+p/aT66Gy0oWbP
IqYbqbs1eBteSQWjDfdEqJPOscxcgcFuyhuJQwyE3HiTm1UyFJ8sQKxWrxsFAMgC
qWTAxkDW7lnWhwPdhvuKBViyZeIV3JJvXkj358EKDv7g4CF8aQZO3yLPm6sv0qBD
MKqxwoq36KijUxdaJbO8h/mB57mgicTtfpS6fhqbqA1DnaK96itcLGXacy4s/7iV
1xeV+Vp8AVglGRt+OObkepj0UJ8qMD2WQpd/07nv1Whas16Ysha7hbUIvShGR8AB
qbUOlTaAtCzVODPwpStrDEHRxjAmAsaYaJMJdTOp0T6D/7cgZJpO7IUobjceo6GR
MCT+nn+DaHBYuqqQaCcY4fxGsvh2uQeTmDwTlpeYiq1eCaD+5crMiPZvm18w25y+
ByojiufWUqr/m1N6Ev+3/wGNvueht84QtgoXNDj2H9CTfQZFe6Smjty326KQpUHa
m6PUf9PdPH5oLIL7zBUt/p3Q/67XVFckZyejJn3C0KvE+ej0V3vb6Cpa4QL3u16J
6Or2rHimTeAhPqxN7Chg7Xru+Gjdq/tPH24wW9E5EwThCsJg+RrSd1YGY7Vsz9Pz
zExjW27y+iikCDpx/XSmuv+2CXIRzPB+Yv9J3hqxjwzsGUBLYd6zLRLdKUsQcW6d
3rzDXoHAkWAvKE5Ywf1CBcbKqALJQ1EIQjVJAAnb6D6kUc/3Dryzp+iqPGedyFra
RnrH2AvtxYc6cqiiOdG8qkQfAMXCHOqCcdDo5YGqYPHugffv8DDYJcDmjn3+nbET
xDehAEynGVf3dXTgS+AS4pgq/SGXNjOPonvGhBP0Sh9gdbEE8QA2QgsxrUbPF2Rl
KakHwCH8hw2IRZt3mr1tUsYtS4V8XQ2apUhMSudN6NmnMQzKQpRvbSWP/7NsIIEl
TuH7H+QbC7Wvm9TFDYqW5K72Bs9bvtaGTB/kefH3SoCkz4FGVuSG+HFFtpNnX1M8
hRAB+iZ7S3gare62qVLeg76/drEoc6RAA8DB7gzlKAs3sVXJkHKEtpc95QKAhyJ7
ahOZ1EqvOtooZ1i/Zw5f13QUlQ6RpabsM+DL+cGfmEvNQ1fs00smOzKi37fg2xUt
Srwk71zO5pAuGR6TFBhH/z+gkrYquMd/OykNfV8RFrzRzUa4WNTaXw5+pgYVoLXT
IBuYRT7CW5/BpFe1lPk17LqrDk//YjWptQ+RMGrSI4WhZTBkLpP1v+pjL8n42r2X
0Qj+EEovoewnP9Ov9dLjoAe49sFLzHW9TRrEVDVumuFZ0FyhCMZOmXoerbNY2CeI
V6l24UTQ6PhmXgOtef5oP9XQ0onUq9y+m8gqOJmCDEBqCqAio0hYsQRxZn/UCq/r
EBQ31ndfdCkhfoAhTrWAMe80w3Ru8SlfJhKUBfLeq/ECiOG8vogUYuQ+DMedD2oq
8sLtIikdCgU1n24p3uCuki65GZDCOn17UKAtBor9yLBqx3tcCoddJM/6OGM2bAEt
o7a6R8tawFfKzQEOplqgqFmxaJDYEO4weUXdPKEBs/wVDArAOuI1406WW7zukmyq
mvVIjgbDPfT+9qyhoqJsQ+pisjlsELjHeY1xbHu+zMyekx7OWA53o8BHWHxQz18K
jqS3pvG7am93KMbyBhW7lgpBICI6zitNJL1dXrnh2Q7YltHjxSg2ykeH8XF4q8FS
x+xPqUPlKEXWl8gCKQgvhSPlm77HCG4K9G/NQ6NjzQiGSD14udWlrH5fNJ2c+Lu+
kA/FjFVaWH78ueQMztfOcv5dnYzEcdsvVOwwfeLvWxJIJTiMRFumhzJ1Zu5dXGpW
QHo9+2HbHUOJMSAPU64dfYV+1UzXIm+ae/qtXkiNusWxDeiMOYGsAU4UHYB4WxHw
CSkpnx0eUYKlgpYL2R7yhC8o68LBBoTxkv9RvvI+t5XOUErhfKCOucgo9yZQR9NQ
dNLebTRwWTPeCiUUg2keNJHux6QEVLMWFXf+pNCJu3aM1TEs/eK1v9JK/1wgsgAq
4CijlKORJ0YAI70IC5f/V1VPCdieXOKHHEMD2vUGO0L77zXX6FZhYh8GbNbGCVI2
9Xmr4GJIZfWn8OJmoA6s6jo5Ce0RcwKlC3PcxaRqSx+B6psz5ArsGRPkQZQ/aJ01
UU9Lng74ACOvj8i5M44K16DA1xKja8FlO401WoI6x174jdJ5p5rGy+AvGPhEwJvZ
dgjMNPEq6jt0QjJH58+Gu0jTCb8sB7BksGD/Z8BcToMH6oU+p8m2dqRhxR3cmOgo
7iAjJBaSacfTYCeGLujTRxbAxFigEaWlf8IA+7A0jLDnhpd7n4j6Vow9FdOVfmHC
QLZVj4eZdHj8zDwbnpq4uKd/uhBs0ZUcdpcihNBTKs3g731ysPp4+S9nULVdL6uY
a/6Ue148ULKZ7dTVp3wiId5raNP5z93hN+ZyZnGT6HqdeWJgKEesWLDWSKDEzvXJ
zt2wTC3RGUdbG/EvwUtOJqP6K0jh/aNipl5EWfTMfYvzvqC3LZnSsSnZAOUrGrTr
sM9KTze2sY5HdgCPXb3OOZu6WDS5Tz4z1QT9hVi9oJqSonQ1t38u0q5Ny4v3zCv6
UhFLlMlVkBJirk7J3lAw8QQwHp2fBkYiT8n53nL9sOPitdxhMpOYvQmQk8nA7Z2h
yXSsVD+q+OVnrKXleyvuDJ2SO6w7BZtXOcYY1d1sFilhikZD87LsxQUbTGFy9xMx
wJNivZjyy3SmjpEgwvx1V1wS+ga4efk/SaLb1h6CpC2y/0TIJHXVGdhowJSVuWEM
8XF72eTAUvgyUcW06fHLxK635QLo3u8FctHzRqUtpsmHrsacExWbRzIGAZC4TVuV
xdU/BTLhTV6m4vvViSCTxcHllv2I0d7cBza1w1jUiAYlFeMPoC7w2O2a6Txy6i/Y
EtANWHhg7StQWDAIWEcvVHUE5VLaco9xZhzyAPjUH3fYy+/SClBVIPUMxKyi1Py8
Bbx5TD4EzyzzGQrOiuzGSW2pDrvM4HTp9x+IKAlcbFJQPPdWACmCjddhcHe+LrnD
zDTNsgRBI6MFr42Gimsu0dvjONZEhwbWnH8WMOfABu4vN+P9S5HuqZ+tp1JbuZnp
2++PE6HkB7FCCfNvZwO4+/Jd/UbV8la1InPLKREL09eCs8hlDBd2HBSMHzzVx9PF
sOYXnWivSpzUCkaPxF6zQVk/vVwkXT7DZ3KAadURiWxm7UEPGQQx4A/YBP+DCtsE
uf6PqOT0SqSu1jgAFyJs4q23rGDLl41OKBxC/s44HLoD9RS6kQzX+Wq/AMC2yfdO
rMlrZShgRHGdZpx+d5r2tN6B/zDoBJ6JvDVS8uqPigZ4Nzfy5zn49LYmtRqkp3Wz
N3oyMXqbwnt/AtGMRoRx1I4FiapckSpkjcJE/j4QoFrB6sAR0esAbqpX0iXjVVet
VZaDNIukRWVFkM3Msrr/rVy6ztJGEQoxhdGcPYXFN9nK2jQZ/HNevNaGzZOurnWf
c2IEzTvIVj687d8MwWMIZfDLpSaJt/Z2a5+RLvjf2069z1bOzi7Nr4hiJV96/jEo
L3PX3UH5vWsVvaDajoFq/NQ8A4TRFD6OXyVrbsfiJ6R8ClDMguumMZCHd9TMMw3l
40hIrQujLbNockxqDFKyUqSsT/1HljuQVA9Xcu2+W4CzWJx9EbGF1St7rRHCSzIc
ijvjgXP7h8NEb0LWRyVX9soLQpVomOCI0EcwtycX/SWiaC7ULdm/9sXK6kIXwEtC
YNWFZEzCZk3gAv/4myRK3SBCLzVDPTt9DhIGL2UYHeXpPIn8YD9KJZ02USueKpft
gb5riB5pnKIB2/1uj4KP0HUv5xcOQRm/LHSxq6muDg2IsQk9TQTBbpNfD54qKOcg
phRN7JrScEpUrMe1FD+XQgzYLZa4ETTkWZJLUEYuyI+NOzs4ei4p0n+A/xP79zlg
cyUuNbblw8srqPpVHnrYP7DZNJjPOWlUK8xe148AUehxhFpnOo8IDQK94gVkPaaT
kxZbIcjNskDlacM9Ne9GvjMyGv2X4Rv0kQ9XCEXAezY49jNgm0eTIbl81bHLGC9G
Fvz4Q2v7YMJtLhaShum+xygYadOoS+sOezXkbEmKaSrBBlUDLPT766TBoPRHZMcJ
+MvmNhB6beWWuys6+AuTXhOYUTQHe35RgTfI/YA/BAUG85/xTTbQYqIGAAlMx2VS
52Cl99x8FxJps482ZpxS+G1yslUOagxTpXPVkaiUKV8U9VRg2Tq9+hLn/aEdOSp8
HFBD43aIuR+Cq9o08Pakg4HblyfMVsAH4FryMNrrWqnQy71nk2R8XyxQTLqwc90I
uiJNnwJkf/QOK56P2e2+ZWy8Iz27Y/wV6hjHYZfHoktF+imb8TFss0ZHLtDzfXKK
3OQf5QZF8EWBNYiJbGe6DLz3l/zZSJXFiUuFvDVZraX/aEj4Z0m3DXrUZVDfM5T3
cmMXVjmqFcGQTbGWh9J6ZUh0iw0vOcOgqQQCpCLeg6jEqJiE9fi85JHOSKEyyhys
LiRQIfShRNRFUL8QXihT2Yu8aEHX5/E4y/KWGyZsvmutczdvlZLPVOW0/2NSzJlV
VqE6vGqda3i7x38IkX6Hwirm5q66HtqD7F/7amL+RvCQ4DhEDJdqrk0XSJJhTXnd
2dRalLkw4ewGyOCGPzhEmgZm9m6ynAeozQvwf6oycRmkb7OKUm0HpWsOUYYL4D6F
SRLJBLpb3c8r1V2njiFNtQ==
`protect end_protected
