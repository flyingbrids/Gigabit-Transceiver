`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
n+gvzq0D2M37FiukzqncbmJTZ2F7mP+Hu/ymY2ocjmnMdb6haqKGVzDXwlgGioxS
V6AN7wNKmXPATSgBVYrhgfgFvHTsYFwWDi3TZFe/5Nws3kztxYA6j2njmnSGFhyA
10aI3gn/okXQ5zDknJ51L5QdWkGFwvy1IOfamItrVGpHl6/+8h2dkKgQ4mmfKEZb
n+LZtOb8Q5tVpt8XgMVohSewVk24U51JPKHKznBMp1VX5MJowIeV/7uplCU5kLTT
4ygiDwzTffT/OyQa05NIPYrPGW9XBTuMHxwqRwxMhBzJT4ijeygVnq42kFLRwU/Z
bNZGJmiT+7onO+tpvxPk1g==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
W+O1BSAzb8uIeawpFUFgiL1cJW2EyqQn7ky0tKhQ2RYqGEgJLgO9frOFSfVr8O5C
ZZInwoyHg8S0JpuN7IybRfA1bjMi7gR5YDU7jo7uGk5L2UG/kVK/WSVtBIHP0QUc
Y3CjenKn01UnaGhUHdzegCRlXw7gADKopwyPsJCNlEo=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`protect data_block
q9X3upH+A9NoIhY4w4mlT81MZpQKLzKN9bNYDU8ALH7bmU3rCBRhLGtLCQxHy/bM
yvDdrr/UUjpI5U0BlWnfllvmYcy8vTTBFv++mThikcot1YHTah4ICY0r0tn+QdR+
nLdo8eJvOl5wlMgI4ID4uiD6YK9TlC85NGg9JmosHNcK28fcTIFlqE+2aYiYjwvt
a0sA+XzCwcck/nvnKYjDuaMsd83RpsRz3ZNEz+LIaz9zH3qvQDGH6HQ18wbnk7zw
g3ECO0nSx0c0EMN67b8H61LfXpS4qGnkKqcnrOhSYDoq+qNL8Ax764JOR5vf7upU
Vz0Vmpm0iU/0OeeDyx4JUGMAmCpEvCVsZfgUMR/Zb90pIqE023mEVnwUYKMReW4U
vRNIff4AV7FagYUVxP2vdumBo2+1QygfS+pgusOevmuffYkgLIja0qoSchwtMItR
rWXck9L2eeItsjMWwNYxTrLEZ3+3JM9jcTWxzLQwectiRQEMnO3XZUTREFsT9z4O
yHLaALc4ys4An+2TLYIz+HSHjYYJcGZnjAhsbedmdfqkl9VyBopXurPz6CcKzRbe
ybBC1GjOiPrcy8QAToJqQozDZ5hmOkWbNAypblwY4c5jgciRyBa5MsDBvJK383Wg
mQISDiG64l1cAT5c8vfvpVkOPqyoFe1xYjNUltNoW17nVrR9esRdWCv+Ye7hR4T2
OsAfl20bhgZ+bNaJ2TsBhbaU2uDSS4MkgyrqD5yCjMY8sJyDxdlvrtyw+BZb3E4Y
d83y901mDfEiarnmNAwmwcTw7zwotCd9iC9tm7ZW2zxNNv083Xe2BTgfOOj2LEYa
PIGyQQsTyRjJFahgbZK2jLWjwB1K4M8jXDDYxFDhmbKd+eYG4iNOBqSiBZx7e8aR
FHYdtLsP6hqeig/OmIFZWn8hezcDzp6F9ZD4a9zSoN9vvG0sZyqw2DWPcPZM1Y4K
Mk6ZBaSiPrMm4hOc/Quu+a+G51um4TTUVj23HqFr9hOWuwsGjdNfkMDb05nisOzL
KfUOJ3DCa3ASIlcRxd28dFr88z1VM/xdvhlVaWwKFxO6DVNcF+PkGOmv2sgtFSLA
4it57RfJdUGJ/5+dV6TKP7a1PsFNEYHw4e2RJNVKityeVh9F08rwTE49hI/QyOPp
21JF6mBNvVHJ7IK++A3Ou9Djmd6bFkNJdqQnG/znxSZxA3IB2ysOAEGkpiTsj9M5
KADkLe3QJfVf29GQryDCf3xAlscr0JbIZQuCqrwgah/iFWG1Q5kLmJTX+jEH1LU9
j/s7F4nD95OWqFFvpZFlWFpefrrEaV2D90m7DVZqkU6OMB50H4CjbpyirOeO+oqh
ljT3V/ksZuD6XubbWb6HRM6uge15qad4kYgfdgbwR5L2nTWBb/1QSUTDq+JmGDne
SEYi/5obqyyg1kpIDdaG9dAoDVR8bgc9mwsFpbYb85X0tB4tE9UMdHxvC4TMlb5U
Bj27kFbLudgpp2N27BSHgODVZUvfGps2gNjAtGb8SfrlOK5wQ9Vp5HpOb8qZeK7n
z+dHKMSspRruZTDrTYrm7rfCB3tXv5eRImhHAdjH2V5RX+IPzQSPogHy0jni2mFV
B3B1gSUraNI/K9QoKWECY/dPnUpo8Wkw/mdJSVHd6W+ReOcxWXQMuMFrEI7L1Ynv
P4zAnRBlB/+hdoY5fhs8ZI0kD9MUusqbGScGaiiF9ETWUWo5PP/8rjAjN1GHxCpz
Zb2Is+QWeQV08P8h9C8JwDchxEnbJ+ywOXbghU7cb0DSAOJuuEiW/ytuRgfw4bPJ
AEouInEMWInWPoqAsuiLg8u/mKRNbQagKekBfcY/k7OYh/7xtHhkdAUXpnQsI6lD
Xuocs+NeuaFkYN/vvyrxc/K3JYT57BLULS+ElUlUuxGEexabtGGwRAPc6/Edvuv9
/2s3ZntomzI+laZL5DuVOJ1Uoef13Z3DRPxSiT2KZ9gJvYnApCNBOGtkcixLQuJp
TAXGFxQG3GCSe2GhRqt3IGWqiOwep2lISjRNoYn5Z7PgxIecv3Yf+Zkm2u01ub0O
FJ+Nw17FgO29h1BNp0j0p7E00l1A+DVfMJBi2HzK6DLrMER+b0by6+9bfB4ypvP5
LyT+M2NUN4VRsq2fkejxf1JOnAHdkdAwgUknvuQVmVhs0AdXv6HW61DkwGZduT4M
/hfWsne87FnzzIBy4OIfq6xHrkuOtHUxOio0YXeYuHnGTSICscWEY8D/qo//USLY
bNOBphVDjZgy55VP6RF3OiDzodDg+bvfcM7QL0/W4QC+toZGYEnR/dy3aGDH4mNb
1jY+tMtbdQ5kNc6rQ2r68pxApPinbDWsS0Jhto4YSg1Hy5C9ZgxJauJMsK0leCwl
FhBI7PwfreEdMOaHLQVI9xHF44Sf+OKPe0NDuxA8ZpU3cTE48qTH7LSIMDIS03zN
7lJNWx+VOHfn8gre820MW53HE882wk6JryY1qas1jj3WHU0AVT3JQGy1CahtAf3o
OaM3dXXXgRnqgTew5UyuWw3mlL5xSRO1vDJ/rDFrUcs16v03klWLKvvYZGekqp/E
sWy5rvfDGSLLeyKjnfgW2j5bVkhVsLHEe8hJboWTDCnWbd9xddkYI3O+tBszOiOr
SGKpAsuwIJ2g8eM5WfyIN9bAMGtaJhQC43kQqgLvaUBr0AXZrt0+tSJRqV6wI8aK
dRgWyNl9no3XiltlnjYRm9mV3S7D73LYN23F4KUf/+2TwUKZW54X2ok7MZsv3MS8
GRRDussD2Se0nFhiOKfUYnEBz6NpF5/e3BAORGhrKlr6Cb9AxuBPlqN2ljbPwfP9
cD5VwzUq12qC4Oe4zLT0JwzrkPmaFB5Gnl42utq3Axv62X9NoQVN9xzHKsvcqFuf
j5xapUtNGWzZ/9CPqfSIUvJupIzzItAok7GttjOKXi5/rdb2Jhu5MF+jf0e+jbKu
vcCWjZ9hIMod2ym25xURe7hYG8SjHVsVqPwoX4PWRWPy18KTb0JeO3ektYlzJSbN
6H4H/IUpWB9f/pfeKxeatRgltOQZvzNgyJndOOMLho4HLdXsHu1S58ukJpQzrXZ0
7qSnvDGuk+pUGgPEcLzhPcmASvG0PnIqOKHETWSBIj3jdGsx1wBcvs52aSc2whVs
NljQSrOhVAYy4IKCXfscwiXEHAYvfFPMWxHcZwblFlQgtlAtRUo0Rx2syiem3UNG
H0i9Vxu6DPEjduzNhz4l6gmVIF6d8G2KM8Dj26U+ly0o1uP/SdgiYTmdzD4kVhLr
4jJqvMZvylaLBsAfHXftlJui73VAs5DNycNunClel/XHex4q2mWJv4MUfODdox8e
b90p8fwzcmfFhbEodHnRRzGjEhJoHXdxlVfMufyluMHiFCPGD0g/JTGEtEXk72pP
bAp2Qclm6gXzXDhAM9MB6qa9FdxEJUvY9wPKlOp6fEk8227sOBf/mx6RWL8MRu+b
vTj4ACZLqwOgwwbeUWgm6koI/jgLMo/wDMAQVYTNKNnyMJmDRGFLbFlCizf/xtrZ
9KIdDz+kJyD+8MupBB+bglwNEW9D/0f7MRVNBrCM88sphLK7gJTW5Ui+J8zQK7+w
3R8sdSewbTzeqk0B9xaNBUMbeqPxHm//DvHE+5Pv05BehlVriuNVuJSbshJ3AZwy
nHC8YMcSVBgLS3eLh6d8xrmyLePXpyd2ad/rXDMaAHbSJDxwZW815yRIpiBJ2mWh
X+z2Pw/LB08LbhZbDBFxLRmE6Yvf0zHqR0J5KXQ63Bgn56lPg+EuVTAz275UOWMR
KZ+atvWdUGP6htqluzD+E5VAfW8JlxDqbJg+DO9NBWs=
`protect end_protected
