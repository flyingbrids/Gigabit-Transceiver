`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
xS3tdeRUmKTVK55xRBQQ67L4XsWAcZEGqcq7bf35+ADXNs1TimfPmNRB0LuCbkXU
pg8d0jERNb2KCKn2xSjf+9SEvWp//zRpbbmqEGetIt7bfWyhW2A5q7v+ZpiMBbbN
72GPh6gGkE5RZR/eNjzzKkkUvOYM1/K3257L+ijzfrFS42SaCNJwie8t6kcne72B
Cc/u2bhbcGmUZKjYPwS1yrYLdR3/6yhMA5qvnAy+Sifbi8K8F6AkKBt+pqngdhhL
ptzg3PkHb2DUqjUKNFvfkvA914mnFkA793u9CfZyVFJtY/Np3cYDWfu8mP3k/iSa
iOwlPz3LNEZKPNRoL1JkcA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
prKfoY/0q/vV76DrexAI1kOlOZUduXtNX76ulgZDbKz41xGkU2EKPLKDENskW8S7
zc/cvvQdTpCssHaR2Vmgi2QUQS9IxyrbgmletcfdS8XHKhKOpuizp3Q4RH25t+A9
BFU3HA4LTVCcVQhFo6Dpeuk7uqYJlXlFgPX50TK0RYk=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2160 )
`protect data_block
iE90KUjt7tWTWvm1B6dGHN36Dsjkd+RUMZoMaFSZGnlNbSKbxt9pfSOck4EfTorR
Q0HeXHfSMCWU479Vu1HZ3dIuVh0cbno35m1V/8MLzSoudpEcd5W97uw3t5MGXG/e
XaDIfp8VKOy+HcP/A5SbCMAAUo59rkKaOSg5mvQ+Jzw+7lbZQeHm6oR99YC5uqK/
kGCHVVfdRGGLyeGb8p8AXsNYNyRztOrs544AqFtWJho5nYngPeAqaaIWf+30rFMd
kSWr+7fTREULmaDl3vgB+PNoEA2B1ojNz29LZGbEjwau1sHDsVgn/BigPPdBlQiY
dTXkJf89YSIKQeC6MU0g7cyCFHEjKF/IbgMxgL5ySSZPc3KeRO16q61jHs9KgKkG
3T+BER4RP8dDbETO3l7oips2ZpTcLHSslh7CktGctFRyrcOVKqFWz0fjZq6y+rNs
+lrpGxKp3dtCbk5bRe2I4GSY5PIFgjqc9t7es0+FBAxLDLxfBBJ7/cfUvArr39jt
us7jWtlaxypInPiA7KJfB3RGfnMGbSUYDcWkAqxYtCSEqiTQDb9HLTCgk8kCWnng
ahP3gTm1Oc7Q+ENPYtdFLZOjCoarxtCfy2sLzXQnJaGIn6IunfEMKUTmg10Kxz8r
MbQmC4l1a1BAm1JfbvrWikg/6ZSuMZ31el1KNj32uP1Y3T7Y5Ait1NBY0cdGP9J1
iym6FxthIYu83xONXnMW1S6Rn3RVlCVYPS0Xggx4aC8C5qeO0gEGlt9Lnx+5bBfg
ql5NsfUGpfPMvwkioR5zfjS4r09EN0JDfcY+3Bcci2Nwj6TCfBgNuI9qNo6ORsS0
icbprBBfeLX/AJWtcCTUilm+jwTcEY2pGAIJDDk4gbUAzL4yzavED2xeOl4rYyAs
rPlAo43pqEFJk1peCp/OwmyQUVRFP4lJmKx/jwgmA5A3wbJBPHFRfh2PDp86QrWr
1AVvCfP7h7RAs6f5dvBE3jcak1tGV1+kZRcO+J5SsLuEYfkU6sQRLx7UswUaYuhA
WxhLql9uPn1dj7TZ++jcaJpnHrBIp3jins/s+1dycRzFVraRFv8FbhcgQ4QWXVMl
rXhJQJzL2kEjuRqe7Gsbqzr442gUG5EF8UT8btMshZYahyeX4gXRE/19lB1DfZfe
ZVysfq0TPHeKWqvPfYUMscFISKBGNFEz+w+IZPtqQiR9e+foX0GENlcvnpXxhBHM
QwXcMxB73bHFqJ2Xdi34frJfz1ZSQ50OuOtyyvCqEVP5/wnhb1T9hvh0qjeWLJNk
NoJ/hRA1/QS5JJ6rnQdrBXTgYvCzMDkkb0U5UGXUFrGOECREkvOxbBFwoglx2WaF
allcOcT8aoHTgl9HzRcS4kOoSeXuWSLA40sM21YrmqMzKcsH8Otp6tOIt0M2WwNo
Ikcah1dMT8RjLhbZrAVln0Tqf7li3lps5y1JgTfNqbqQ6TojG0a2pUOKcEbGAIKJ
ekac2BCzVjSE1CGK8Mm7v/e2bByuir4tIREGbtnd9EsmRTX2e0UJBL3Z00m4TYER
OoRUNv6Oqha88X6/kuVcKR1L/VA3Nn+/SduHBXNeHZ9HRD/FsIOf50UMtBLBWvzL
GVH4Rm+7MH30eY1j/7i0Txe5SNGqniK5nUEQBFqXxKvS0bIF0CAUsIPBKKWBbcX6
aGzLwiQtXiQgq3MJDdysy8B/2sDX3WPaj0k//q1V1pheCyE76jLvEO/TB/+QMMhW
XVmZxdy61Jth+D3m+/7r9lyBoKIlchyXDsrMkKHRVZDFw6czdu02JJFxmnEfBvrQ
Hu34GkdAXDL0aBM3+PUwUuB5/KGDaJehoHZYEzETjUDtRwlL2j4M50PAQQ53JRu3
MYzUFrjm1v2yIxvS5ebe7rFuHskGkvHoyx/b6TWLfRqnlpi74fZp7UBo2AE1a70f
CqBHOoeIVBgPZJD4n+3WlXQjCr5a6I1/dRx5G1lqLntBSgVvq/rp9rfJ1jJoDFCx
6K+tUX3X82TTUUU1xXEeUXVrXkaxgTi4n63tmMDkPhxlZzanNFXSrJxm//xypJKl
xhgFim+OkpPiCs4r0lMFzWFbnwvrpKAe8Mssg5kBlV7Xuv9gMh8fL/ptJqESmJKL
fcfSLug5ZjWWFKIdAEwRBYzoazxVEtneNvfhW/t4DxIFnEBh9+wLd0zz5ukjm1vn
7/4Ixsqn+MEv4O3rHovO4mg6eLgpCo18TTnFZUmYO+AEDNtd5bI/IOV2WcoI4V3Z
qBBE6kK/ym5EjHNwK4PMOo/QkQcqC7m8B+NUEDK90RhoElxbq1yK6u1cJtrHX1eS
X0xW/VUROeXi96lGUxlFXI9REyEHzqI52XxKqnt0NakLlNAsxPUIPJIEgT00ofNF
NfjUsyH4AOsVc0P71YVJI0D/3R1muVjLvClE0zmaRo2IIoQyGvKm3Z2l/llw+Bhk
T0by4DOwlegwLwhFbm24pfvErdfrPOu0w2feInWw/AsZuLoExkaCH7HB3PhEX1PC
+M1MpcrT+53J5bAVKDnp2MTxQEqWa4+1ebWO6+BkHBX+1ohcfFDjATAhUwex5GK6
i1TgWzrXm96aMrukLZsRRxQW+A2MCu5AcBH/mj44pZjIwK0pzcYVMLqcy54vgXvA
cGNgFrSo0MJCeZ3kHJBhoOdSGnxg//9hqHHHKJ2eeQrJwmw9NnoBEJ7lNUezX77R
Xh5HAwKTWxPZhrnEc/0FqhAcVovxFY/4ALDvcnX6N1CN3zPkYZE6ONHssvNqbydD
wLcoeapGi1Fr8zpIVbhrTG9N/7pjZ0G4Q+SToL4fQgj7LyYyNxCJz4M1YSG/EgVz
abKL8yaWEFJgUm4S85Dni4MQDxVX7v+/a5OCU3qdAILgxP258FFUl64D2FNtyisn
`protect end_protected
