`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lOMHhhtVlMTV7YvD7KcqOtCth+Buam+AA/vHvX/crjjqFsZDriaqNQ7P4iDLIy5X
VklWXunN5TrPwvU/RQ8XTCcy6HzjEmNSMSnMfHrn3npWc84vf8H7ETCdMqmnUB9f
gZyEjYbXGlHL4xDPQv0Ael3i7tRad/vlMqpAq3gL7E3b+j4QHfASBG/f8EW4uNKq
DounsmJj8vnxszHcAOZsEyEauvcjPqa+fiIqp5GIfeq/uoIHaoihHYg7XNSBEKjj
REpN/ppxqkFErYLsamYwnDBKL91PKmXjTtHY3Cdl2G0VmV/YYoue0373hmSsg2KZ
UPqXdbMCDTJf6vmlLRsaXw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
tGN7l2OWsJGtJOuemdRUlCnDWcK7ROauyEJagG8kjV6DfZrXUkyAD4mFs0CKiwiq
3ngz1p0/9XvZmrFAch6uozCXAgTXbB5VwhBb81L/Kf1I7dRlWkSsFPF8LkJTO3V7
+miLPjkQu0MWzwfm7X3VZMBp+ROTr7P3G8OxF1QNOhQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3888 )
`protect data_block
7miBPwgh+r+PCQ8GBhyTv79uEQ7ffPMpMNRdz6vwfOaBe9hJo8f4HxWEX3bGh9Fr
TzZqaIv0dtsfiPjCwdbHgZ8Vr0MyAHefstUGO3Xwr6ziUml7AU6JvBRWpUKDZb/A
W7GoC1rYQmXAdr85b8FA9kyut3V01ZUQ67TAlPssF4sQhpvJkR7ZK1bbZIeqrqkM
gw6Ve4bLU1nm4lVI3KQZncz3ObvzALT1UJcY5rMKOBPODdr/u6Si62b1ybywHcrG
SiGBt2i5kUodh7n5dM6ABs/QMgokjhZW3esScYiIt8t90fbtPwBMFBwf16XQZETI
okeV27dyek3HCZAFyTm6yz1cAH3PQ0dATYO28pl/GMNadjU9anJM1G4Pmh4GpbB0
5JFCSlcvVSQ7vjBZG6Ecu0pqrgwmaJlEaDVoi1tz5kJRNJVchln+303QMcbkA86G
jrU+ah6+ID/R1fVQohhUFBC+O8UYPA6t2jyrbaF6M+bLsA8FhLkiGhZA3wGGRWG0
li/6xiJniwj2gETw0ElDnc8EfwyPvF6QjfHFQIwJTdpaUi/I1MgsLxPlATZ01AuV
03ZkG0bTYi7neYBMdzch9YZSj9M3smEG1NXYNsqS+IkY8t9Trv3kPlFUyWD5PFCQ
Gg60V3ZK2HbDrZBzhvT/q0DQk/KViuSHEQmqUI+rIwvUiqGD+Spj96M7kohk3Yu6
Vr0RPbkvMOwi+XrMqqoWZJHbCpaawGQxlKM+/ipQ9vwsNxQSw8VgMLLpfuZfoLR2
OxrYV7FDRGarl0/MP3x1lQIbL2toPDpUXiWtozpAkoPTwo1SZXmf+hYNS09rlMMb
LjbkSvkv9ymtUwiDQAISAfiXZTlcr+M5YuMD69Gf68NfOnuL8DFnFh+QmXclL13H
HdPQa3WtgIvtUZtNrMAhkpWKKYh6SxoDFZLnqo07U/OO6F1Hq50xOMOs2vFAFYNj
MoyTDrBtHO46TuBYsBV432twoPYgWf26k3QfT1lVAylRWCU4XeUrpKM/jIbwjDDR
dCt/mxZ6xUsmj7yvOu1RkqqKFUcjsTVbGbFjuMOs13Dz0n0/az12GMWZ3nISXsSG
mHpIilJWWqFVekxevEGk/i9Ep/KgJ+n2Tjcpfha5GcVelkR+jvCcwSVIzbVERz3F
W+CvyP4uM6MUc9vv7fFAM6wX4qPPnWyXySyLpltn7YAZFaNFdvynT8uD0RGxi9Jg
uOykFXHQD87znZaOGaNIo/FJE/IR93yvQTnh1hCf4dzodipbicn/ROVEtQNpGSmZ
khBm/bQCCwn/jaCzS0lXHXOu4mZlROLJ2hktqUb+YDb5C+PRIS+/HzcjurPVTCkE
LFqQoBV2IJAKZPfg+2yZRNQ9k+Ii8y402zmIVmGu/mNQQG6wH+mvNLlKxEUsGq8i
Ym2TFwEDZcNpauTfYHpLfSCZnCeToVyYpS5+mIlI9L52Lor5XXNj3tG5bW2OwOah
AkRf8DRxyNCFv85d5IrSCmxxC/82Hq3kmGkOsIcoMPZbHf0z7o0BfiNC8N5GxVQu
/30zRom3mwSWoEWNuMZ2azLchr1MMN/92TNVH2y5kS0I3ONoNF1403To+u2GP8YI
jvUg30TckCUyevpD7QQ36qo6wDoWCJEnuMPWzsWM3+TkVnUUbz8cQjI9t5dMo4iB
Rt5eO70iBFLkcBvdLONatBy+t6FbKsWUQawL2Ub2QmO+uGfh+abFxTeYbht/pLBN
asgRzTXEe81cvEnbGwEDBdJhyYCgYcpaQFFI+2Df/9Lkq63IYrqig3+q+L46TaNF
i90CC4uEE3NdorrMoMN5KcAnCEEm8IFj1LWPkJF1894DoCj1lG94C8KzutzrJF0N
LdwrxVwVU0Mk6/8GKshZ5s5MLH/oPlAcSPnYDMJ4phcTkehVEml0QT4MEmZuVUT0
QiRp+yVKQk+9WxeHRmhXXxheGYW0Z6pB/3gYtopAKrO5vkWzZPd9kPQEI/qaeCia
hVerCvnmt1Lco+8oyusdq+Wmx7JtwJi/hpJn6P0h/uCsVcgiGeiwKmTHVQcvMvcR
BflQHaqsbvNGstFWAgDRcT0byPl4BgoKDoVqeNPkBqHumqxCVMwjtMSy0LL69V9c
jI66bj7BYLHE4i6TW6myEVE5umqq0rVvFBEkueHIK3FRMwU/RLyB7TJwzHs3NSKp
IUPFoRddtAjXkjcveph8qx4Cr3nG/mBwIabDvBG4wQ8///eesjZq24RfFmgGg2pe
5gJ/EEGeZORC5QMwR5/HIoDnjBPOJ69/vgrq/Ok2wfdgC9jCjkpZCTrxCeadeu2y
d1aBO+/Bhjk4/RJrycvRpZsxbNzazXTo8pe2obRFWBmXvVvUwTZmJ0iV/dtuLnAg
Hml5xsrBUEt8noTIiLtr2D+nHmH0KEOggr0jDh8tKdFzxZZYmj0vBtz4/8F3Fty3
zLYcIrWullxd8zMe2mNPVIJiuzUuZkwkQoTEw72Tf14uivFHlTgQYL3/BImkzQz1
msIcF0zA4KEm3qavGhpdmKvxnIsjXh8B6MuzxTuBka/BsXcAaV3UiBFnIC5DAAj7
DxniDUKXZXMpm5WUZQW7KqAPxUq1Hlu2QvAHXbxUv8TOmrytKEtO0XwfzLKUKjZF
87NBa2h8lOvS6HqzVHYz4bnVIH0VVz2JESrM7eoh2FViq7ccFARFH3zJZqklgWq5
OPCS0In2haFs4c4hOAR1qZlLZNDECswOQqNyaBHw4v66yfU/eMwkTe5+IHnQeiA+
ssjfoGJQM4x3aHUwSRjr3U6Mg6XsCbKcDhOHEixrZn6IG05z8L1OtZ/M1fCdyvhh
kqDWj7CAi04Jg4F4z+9QA6Ix1QphXUkRd7/9FjQJ0ZxkoPsi1LZxUskLQpgx4SZn
PsTrfojjVYn9JNycufkJ/fwK8NuYUoA+3eAPonSmlTn+u16/PqibHpqIiFyRTJnD
gxcIrYkPKjBR9kd9YaRfz2vygsPx1vYc6KiinJZvoDFGb5DYp8+mS2i1LJZ3jyb9
hlSOEVwEdtl+nBzUx0T7Rwy/1n4nsZv11aZ4cVKM2CCO/aQRaRSP2TiCEB03y2tU
ucvLllMNhlrsgmD6kj33nWHaRTXZJR3/t1DrFbP4BF6QKhe05AGAoye/NAkEY4D7
Lf58D3PaXIw8qAyd1p6heGSN5J4+XsjTamaKJeQU6Xd/IgW/WuPhstqsKrQxnBTP
KTWVoXQ/oWBIpcbzkLuZ+XnuZpVSd39cKs/0gokZWAYjohKEyNSg2rSFUV90gTjJ
B8BHM2XUIddhOVA+I3VWhFn3fBy+OYPbgV6icMhan+Rx/Jhs31vfvzQRKAMIP1yl
rhii1OzMwA6qNgEnlQXw1gy2gHNEZdsayKiXRfLmLtLOfonYLcuuPrapZoYVDePL
ydWr+GbAKH+WwlN13XfbTigLfIHfLfedjI52KDD2ylzhWSFuVNAaIN58/2ADL/fc
bt5orh5RxZBqIjUjRc3sMCOTz4MZpPWwG5bb3ZeAUjdxAtD25zdGs0AM12xh0wUy
KUCdE8dr4YUY+pjf1ZibZdarZwHpcFG6stgOEGOYg8PjPKbL21XADue8vkyuFx5j
JFFHIUc3k+fAzjBmnLl8Vk8WBl2cCDMMkDg8wuQCPtCntQN++IG1y+EtNL+1CKmO
02KS1UUCvxGU3xtLcek3H/5DYjteQxQlpPYShGTLVTpiY3Nfw3VXOCQaxhWJ/ib7
z+IIQKen/I7uM6hG97FBU0eoR44EnmbviB6Wr4hIjy0K+WLkZvO9aZ/er10ZTVv0
VzmRt6lghjl7sUD4RePC/vYn09hf85K+oen+FZ2x0AvmucerU/CcKwBKrRuWleWN
VY1MwBnORdELoEeRN8MNtufHzgyYqH4yGVKBMWGa8LyehoBV+j7FWjsRV+3TKZ5E
5VPrIHhOBwiSaf94EkbhaI3v0Jjk1aMIM9NDYf2Qw/VqFlMOI9nOPZ1VhuuhKQ5V
c/9D8/+HyHHzHMgH9OmQb6Bv8rw/FyYnJnfuM7lDfEYCSi+x4fMSJnfKQOZ7K24/
eN1z0JSXdMexoV0fVCMegPQohU6/V7MxENwBWfUHx/ow5dtUh8xk3gJ+T9jgL3G3
MIc/1hArEczU0BvcNnmmCHqXC7TSTSTQOeKQF98nBtNekWf2tIfSSAeelvSOhu8U
63gfH27d8AtA9Mej+PPKGiw94ILlB/eD/mJ9jMXMAgROqIgktJx1pIHkf+LMYQgo
O/yteREw+NoXDEZY0uhqYdL1cgLJwksZB2O0ZtzsEOh4bu2eoF79mrEgguiQvStX
Nn8gEDATDUTHTDyEa3yCPOHQPy+Adj7Wj9dJt028lgtM1a1T6B8ArCSW9XcZIhPK
CxkYntLbBtW3zGoNHSkLI6dsSsx2xaQHRG+d/aYIqVqFb1GpFxvyW8lWo10dJApu
g5gzrW+9eqvIfFcsqYOFnhHoh9vDm91PwgSvZcFT51RdAhDggipY0/0gV21N4YzZ
L9ANsjJqeyLSHnVcF5nSTqtYfgXOhp+CefG4qr1ibBMLRKMVKv0YP3bqjDJgukcz
l5wPyMgzbLRhVncG4W0JUq+KRENh5LqiqLegvwS0DjQ4HKGGdGBQBPFyfK2CCO3W
jG7YGseMr9FEUWWywjK7qFUMR9PgPCqknWJiX2sZN2MgDmuvMSm/x5rQgu4JVzrq
cmyuTfkMuW3jy9lADk1tnmzdUXlNqcwW027rbOP5aUPLqlaLmcpVdnoueHkeRJIq
bMkbXFpvZK+gbJ6a9uc2ULuS8HlvN0VuxCFIKR7jETeAhsasNpCubK8l7J+8WrYQ
3nzUEu/jomxBixt44g+5feTTdby7SW2Y0DX0iFjAZhB/D4cAtbikgYBpHw83kFL9
YTXs6j254To8GGl4It03PQ4MAK/Myd21c8ot1ZjkzxxFDdc/yU/naTtCuvl9ctzq
FYun++9Ep+OoMESh3p3BXcrYoFKph2qBBjBdMqbi0x8Rk/ecZBr+wlm0hVMkaEEd
c0PpbT1IQRP8hnO2P0oeQ9HXoCVZxdTtL4yu0PDjdmotHbTYOB+UjpAxoIgA2EXm
/7fOvg6cX6V915Jtw3yubbtYnFd32xO7kmO8GJ9kLsMc0OsvTMOs7ueVSQHTwuSb
AVrFSew2hmgd3b1jLG/CGzg3+4XX+V77N9t8SUh5OvChN9OUg3Teo0ZYJJk7748U
`protect end_protected
