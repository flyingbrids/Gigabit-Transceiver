`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
XQ41xbr72SbyjdkZiWykrhih08JIW+fBbGZ+SrQxvCwqbQe30ewISM5Py2RRHdv6
P4GWsqIt7uFf8b1FvWwp8JHS5YjN8NolNcJnJVMiNsO4WucVDvUGBZvlMWhY78fF
RdiK0qK5NBH05+6NLNMkY16SM5uxLAjK5c+HfvCvitff8TcL7XOs0pDhoUFaZsId
wSCIqXSoeytunxGFaiqRtiScnZwKvaJHdo65UumrEjPobr7Lu2iXcB9a6VQtaRfN
VuJNFADZ4BYyggYjdOmc5lgzF7rmvd3ryA8LNsTxyuXANL2zCgBDWTMZJ1xsgFnT
Lcf2IZjfPrK1DrZUE31nyw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Ud+P76NbpVVA1EeP/gkUTKay77Wqk6juFUAddny+54ilaqjHmO/CoYDT9MTsVPZe
/IRt/MqvgJUyvkWWzeGebA3iMx0TdnRf35v8hnKAPv1vNkM3w+JoNqkNxGgy3lYe
VFVL8Mryx4KsCYhBl4CJ2MIBko/11xg8fGUYvCsdXGY=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2368 )
`protect data_block
1p5ji/Inc1O8mx/NfEJgPRyEagoj2e3mu5WVCsLgA9Z23jsc74fQaJC5QVFL2icc
3P3fmusb9Cit2+fGZ+23xhG1cTsAPxN8nv/caJMgHLijfF7MzXy3fhsM4nrNVBzJ
kEYZ0Ng++gSOx2t250TmGOF21Oe0GyIHH5c6dYZN1wqMDF2Q0PRXwaHB9QTEZajO
1ng3y6na98nSxWZMCYYhwECWr7yU4mTVPzgMW7O+bxZSffi+54znxM2bt+AjLnau
lt+nVO2IxgjBlWeGChoRU+UhjWpKkIkQcIamM4UAnqD2odsBb15a6C+EXf51VK7R
mvvwal2rYA4snFOl7lhvkI5IbzCvRMSV14+avBEPoD+piiSMVSEfinRMIjkPO+F/
zmAAGLceM/bD7n8kzC1q+cecDmsy5Zn41ww84eRFhOAgc+7Tl3rYbZ5St2eBUp4M
P6YChjiw5/Rc7YC8cuzwnWM7CrAFszM0WcuGsjr8NpJwI7fDPKKzaCtbha3hIvqi
k4Qhe4rbvyrSlcXgo6CBM7PYAQ6RxS+u4VjLOCvKKY/Cbh64Us7EV/3+OEpbEGKN
Pdxy3VmnWNSYNWzH1OnCzRh+5gpllPlszpcNmUd0fXjN5qQ4rmknY3h0YlFRa5Ao
SuFo1Q3qAtm3lpSnKfzm85aqrL/Jlg+A/PPS9S7Vc2oX4UklopI4fH7LGkzg7BYX
H02QeXx7IOX5eEeYgQVT2hALJ542UHvmsEI6rBn6bAm8w3giebdgNwjR7hgVjVbg
m8rClmENpIcxFhMwafXfoTf5/PSSJ0hr4RmiNig4QTL+HNJxQX1Is6vllPMODVaV
5fm7rI2uPL+EltvVzgvLEkCsQZaf8dT8n9TCTSqMo3GqGSE/KTqzekyRjF26tf/m
yNJ+KYKeFFKQk1pDbA4YPCosOm43f4D0y/QdqXvprsbM4RMEI+d5FZoQvtO1aJtj
P6oUD6dLd93563OUk3wDm0ViWytCWoZw14VV4ioPngXv/n2tEAD6RxxqR8q8m7Fa
mJMJTy9IjaPbsrkXogCyA2Pht3O7IKtiA5B4ANrP+CB872JklE6vzphb67NwiKl8
4gktaR0xLUa6V0kDYrMY/uOUg0O9bHWfiVeQzw74bru4HzYf8KVNXNHZhhxRek2y
XDyWRGiFAEfhT266zOjgOoZQnNLDXtHeqZ1UejbMtTG/MdFr3XCrJVIBP5zld2Yl
D0QcBC2Lkn17qIUrSOjIe7yI11OYghAtmNRkvKM378wZSPCXDD47bkPVmfsXVuHH
Z1npCmYTaEXDQYbltjg4YGuu7khrGgWvf9HnGpvPF19o/Nk3R8Sl7dkatksg55IL
BtnCCxw1uSP3Gsb6k8TT09snc7TNff8AGQ42WEv+ya0mz6Ud2BK6zq+tQfyDUQWI
ejMpzlmsf1ZA1uADJY/0G0FAlSxmSEDXAsse8tIaGS2bc+BxOVTrZMy7pTwhI7of
diGOlLIar6j23WFi9ThPfeJAVYQKHIDd5mxEyhBRL+HEZKB0TqcQ+jDxyqcXN4E2
Ync/nFzHEQEB8MVNdMlGdAx6eSMGf2xiIH5fHeg+ETfFjZz3u9rkg3Qj/DCfTaoN
tE7GQerTzhvgZbqkW99Ig7lfACQNJn6OOQqokSzTR/TqWiJGMJBwlmAH+RmWPToG
kbmp2fIpF49156FrLcvQyr64eVKap/WKysd8AppIP6+5Tm1plhCIwkWujTxcdrEK
KWU+D5iTIPazgEJNsSl9FnmUGhIKrVoj8L4vnXa3zS6P3P/7ECnobZk0VTKaZr8U
YXkQO/CQ2X2K+GZ83V2aLzFlWTxiGZ1nzuZGfZRAw3jjwLgYuMHGnGpLxhu7CY6R
2t6Bkmo8WUkv9FQeP7M/wIPFLNgCovanjOKGwsApH8+D8BwjuNg2ZGWXJcEzeTRU
HpmJWYA2ngL3rWfO4fK6Pu2PYCdMPewHQasssy2K1P5de4MnbaKghDd4tLF1pwhR
/BrV9lb4m6/yp7Zf8JZI7WTvOvqMPraq/cj+23sufflZjS+vNDLQkEQzh1Vn5d6+
PI0sciIzD8HH9v2z1wH7dhSraZGT1/MCLyHoE5Jc91C8+eIEE+jglChph3Jfntz6
dXWVEQUtFd0+2V8dYIhUgMbsYYQMDNvkP6ltOfPSAr4Kf6XvnzKII7Wb9BAnM7GJ
GcDEPOZ6xQDoUtw5Ta6373P13hVuOTdaxrFV4YtfhHCdeLrY/2WljfDv/KMv34Sh
Se1w0uoX5+IpwdM7Zu+xSzOdfHLiE4QWKnfqMBisxIAD72Z0fLS8zyxBLoh9LJSd
PSvUyUlsgHpZaWv5GQM5h/f/N3dmWvFzpvnFC+krU0xWUboXgG+pZEw+QwcE6D48
2qByyQqPQ1X79AreTu2umjJfD0CF8lZnnWCg60bBB+InvcRmOIzdD6ejNu3s+JZZ
D0eGnPxlDdRWiDIQJI10t9yEECDESe7GAnhGSHTV4P0OohjJPJ7s5PXtg+4/4+xW
7qmOM+D1ZMsmmyfbKj/4oz1YoctvGo7X/4Ow5COh8mYzkOWOic9g0Hb7VWWmYWjg
VdZ/CkC62GRsldvSgESHJROS2z3efE/IxZV30egbN9xE6qCLhMRHC7kzajAVvsh7
W0SWNMV6fTA00sQj+pTAO+DFXhoTglBQfjJvpik4ZwDjzPFiI0bYdHOr9lUfSn1Z
FzmwxLxq6h8PcOz0xLu5jCDIOEZK54B4semJCxDzOihiFBEan3U+q8mT74nQhLFV
s9wFHlx7ys9YbACBnWwKeOLpetRCNhUxNqJRxlWfEEZ+apFfwZfDCIOqs6KNZnRx
JNkSCLUglFGs3xuZy/nmx7qHfh2DaajvTS4QFEwrQEpns/R466b8wBPy/9v0tUfH
FWTea0bVxBeDVv7W8QY6iHcrwBK+vnnOcUyr4pe6AgnJdap1ArWFoib25a83K1pk
OnIkWwr2PmEaf84xF/TUk6GlVGdgh5/zBlRTPxndV38emtYduBtk7kXc9gO1qDV6
jXr71i5zo6Bj7Bg5ceLDtRVTnGhJ31FJWaZFnS9UojNimkyswe3r+He4f3uGOUGC
g/NM3Zcvj63vR7yMXYVWOBYuwETovLl5xSgeI/RZz63FlyZhWcw6OBD4NHTOpfdq
D3ej7rVehIm8W5npkD1VLQ==
`protect end_protected
