`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
xOGELUQoZlnPmAQg3c+zx7EoI0hcwxTo/Xy3y+OzpcbJ8OKUENF0fQo4WMP/WIGg
/GojXZVfErHrAlvY0QcipN7yd4FHFRfw7xRmoKHkrpdekKUyskWItwAlL/a53FTD
vIoLuD4NV0iKEvPLh0c8X0apchnV0EbJfNVNZqCmrhLU7fa4YAS5st8Au/Kkg52/
S4xCp1Ei50F1CK7pCPu7NvymLF+slv62fYOaY6jUTlkciLDxSjlXc65urGLaJYjN
feeeoyfL4emUakwAE1mlHJV11x0jT1uchS4E9vB4XOT4wSXexwNtDCOtfuYqSelk
CAqs1kwzGiqExJR8gSLoSA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
tPJQL52fxlOWuNYVi8EvgecAZcrl3I4PzshV0qAJxAq93fS3ByX5p1tQv5DjJ2zS
FapXlf4CE4KdSeYcSbPpEJPOV76UuTeKniq60FmF/BUsLr/z+iY2934xWrJLkvvh
POPsMBQJeFSEfUYHKPUODeQdvxA7yaR/JYjcsoLAwz0=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8896 )
`protect data_block
SBiwgwDpp8EU9pyFpXVLORu+X/ERMLU7mLO232p6IGBFYSeTP6g10K8iA6r0V6ns
SWz5BzG0EZuBnM1EJLm1MtJhyBlyiS4Qy58RM3DFqXVZ3fn6ZdPk1VeFn9OtHccL
mG8rO51J3C2OvGeMyIa6KbACI+2K7EkXVMQGQt8TOAnc3YRiZGmLEPLPgiBL9o+Y
cQlwuQZCHpbmRj1KBkpgOoA9v/m01c8bY1VTVN04N+7gf52hKAd1CVww1C/IlNun
PveHCMqTZqCmX97nasu5vkVhFwOuW7H1mpcFzXUAdmrdNsrIcP3dlX+K4OZ29aXx
N8IH1UWoypo3jliLIX+V1TTKrFWa4tGJsXONBYP0iQ+jlm9hWo4B0x/8IDBBeYw4
lqTE6xVQmLugoU2VHioJUG4gjskgvuPfSLuBlXCLqhhd+iYYRSauRd+A+xdFf8Ws
K00qdxsNA8jZ2tF73vQMUznG/jOA0M+f7eNvH79PRJgvVxc0v7Dom0Nzyg1kIRVS
JfXK3mufJWfzsRQIFVYPpPIY2fXIX4dWUvMTQ3gEIbL+n+eRcuoICL2kZiTy9XPa
lUqFfKiu/+Bc/WZu1/A/k8QyN/tEoD/oF0B84bmF/Sp4z/qZMvVf//PUiewl3CX4
S1WneCsExAV3iK1AZMbbPUdgmRH4X6HOsKw2J0QpPYo31g9b2OG8vNLLLd9i14jl
hfEdRa7Nqi8nDdunN4874vrUntVUre0cSZ4vSSFrv2Qq2Mw7Gzk2ZyIb5n6I1rTF
Qa/FQwQXiIfrKsit5lNz58Af8mrQxMkdXTNNkR/RpISPa8mrDgRZ7YC9tU/tGuJS
WPK4CXZsrRiS40iDTc/RLtyb6RLtiztggCs78z9VCxHyOSmNR2YqhH2HKL4FcLf5
z/gSIdifEGn2e14Q8XrrDcq6fk2vH1YugC7MSxL09nmtM0koWHFXutCWlsC2XLIg
0eY3L48oyFc01BOFNxfwd6cRFUkK6G887EteINcySKwDA+hoK+Xa/+MCJYX8XTO+
xViMVC194NdGmFpq0zAzqkCpkilZIg7cfqeKd2/B3i0sLwxqz1hu8vrEZkHoF6XH
nqEgHkrOklfO+X3IFEwbg9DzEy2O1zD1zhHpVmSi8AzX4qUhjzcpOuD3B0PJ62Ve
VJWqMPQ+qPyqvjR19E7KBYzjKtR6BBQvg213o/tXVaHYATo04FHfvKZYBxBlrZPf
a7K+MLGVAFugxRQllAy+ZaKA/H6gCg7aCV652zYU/6ky68bAH8zKBR1FhIEO3tLn
IgeT6LmM+tNxdwR1m783FCXf8yjcsa6W3ImtQz6fViEzbjQcRdaBTCPTdiBV61xn
uK5/+uLxUMCCmGl6UUGlcfHa8PVuOnf7eDjGFku1sS4VlwUUvkCLf/g5NTFP20KG
MNH/LrvQsQIE8JuXnfVT5aZb4GhV6TwK5BrCvpYdmFdU/WZ9upvvqsxAxHUP++nV
EqQvKqVccPuWxCZjmhyUY2iBrTlZrD76MDaKyM+kFwumw3KIgQuWWvGqh4cLGknr
DySYADm+qLsHJZfOFzGmeAZkoCErVSEEfizstvW1iuS2dFiIYRKhgEh0t1dkdDtM
GtEJNp6BCKT/3N90SPxCahLu2Eqw52wlPbs8NhZCXGdHjpgefRndoT8TJkdomDli
toQ+7wSMxFt1mq3XWGdmAEURCV2mBbQZZ7X7UoKK0dhCLzo1l51zbNFpWJgtKAfq
IMChFFEOSFE0j0tCAPKJUgiNnWqV37rabg8CLfxMfpzJvcQFWb8blDkRRHIBcGY8
ZIIgJ2gjpJ+pN789Y1ov2kbNDsos+9ZxW4Ihb6zNCHay/u/C7+gN64vtVpoqrG04
v+KS4U9/X6iIj/XP3ITQ+akZjWopQdjMAyBwHq3kj8pJ4HbuVNiUH9wyA9yzwF8c
vPULG7wnmwZKfqC9faVaMQlfLOBYQN9L6vt1LZyuF8rs+LYmEYrfp53PLboNNTXx
lYIhjXxAXGcjKLaEh6v5MMyL4wkgaBP6609sGd1C8GhJ+zCLoLYMJaqk7MAt8l5/
G1+h0wmL5NzPssgVoRsuAMvrPrNyNt5AhbDkpG/Ep9GxdQYiMVwc2exWmK3svla7
5TPTqsL/Lg0XryTmJyF9vvNwM1r5jXz8pkCYhslwJPoGK2YBqwu1v56k6H4csOud
rDLBOxcFSmM6oTibV95M3rXyfYIV91zi+P454ub0JVYSo0p4CN6fJ2pm4mS4QriE
YHY5ssqYj5NQ9PKSMwl+XkEA9Oo2BmQawlsvasDhAOAOkFBecDLQIE7baQ2bTMU3
VxnaV5AP54Su8hoPlgZP3eYvBH736CRKW7CMx4xa/kST7XzywOt4Dc01pEnkEdz2
GXYIY13kfpqfiA/TfDZIL34JS8/26oxgNQdBNwcgstFv7ydtHlWYqqS2lKsksRja
S0OYO3zKM5QZnH3oVOhk5sQ6YNw3iEO2DtS1JiAuDBETrEXAEYX84WFSWP7ZxZOR
6mJ7MvMIwWY9QhQ+2eooGbFH0mhVuLVOUrcnhAd+fbY/GtwRroK1OZ2CwhSLHJtt
FECjfA1ae+7UQQ0Bf17SRsSQfyKglnuMQjb3kwqsTLonjL5nk4OJ5gjvE0H2mHfl
2O5hl/jtl7P3bHB22pbEIor9iyjlI2NNBUfWHgce+O0fVbv9lji+OfhQr5/OaLfP
LWttcTVJ3zBYbkiPVvjPu2qzfaeDLpnC8UV/+SZzeSKTvCa3vShKZc1WFTqn5jPY
ArZMmjUtqUStktIf/iutuq83rCh5lzsr5blgF5UmzQVUSlqBNJuKYI1q1vvFkcl6
pIMxxLcUhyY28O9K0n/GfRyDRf8fGDgQS9aLFl1Ns5NIja0Hu0ftlkVL4iX78GGI
5GFIkaHTgPRU91b3leKAzeksGAiYrdO8GU0tBnVfN5XEU5CUVusV6QvT1ivUq7LW
jJrXVtG7K4s/uV+fiG8l72UD/VSnwZb2ZAbIvbJvL3cs0G5f2tkxiIKT4LVvcluC
/D35C63VPPMnyRhLobAlw+U5IpRRwwpPAvbEUcdPar1ergdJTGQR74kExQlNjVcW
01I43XHr3eq9vclMmfS31WY4Q+AngKd8SKpJ0u6Aoe9FyaVPqlZsCUa9q8EI6wz2
sqRQX5VoxZN2gEttRrRxCJXoE5PpdB7yHPpwUCSa+8yBrLmHndWoa8A+3ORnHt3M
xk4rWrOMppasY565XEwFJdkCNwSCiqqzyeMf7O7inrRVU6PSXuA/xeZaNectbOdf
l4nM0CQl1RZQnzI8C1bLrikE4sc7H2yH0lIA4yBqn/2AAFARH9BGrtYVcLOK4kwk
Koo6Ho+uX6djZvZUe5mhgRFabUWexipwUKYk/URUpIZNkmkxDz/Bs1+tKzh8qOoA
GaDS9YKfDUVojKDK9Io3MJtGPFyJcxaf1Fi6Mcgq/VmNLERHqqDjGqRNqsHxH6B1
byC6xjWm3/gPoPAbQXkjDjjdteSibeKG52+iVAnUhWYbbEeQf+1ypVEBll2ymVIy
tPPhqna6Vxud2PmIIDp2Vui2w7WLcVM5DS9whN2jcRKmsVq4rElZPlzB+KY4HCf3
ZnoTTqMYpojbpsbhOJhiM0QWHEx1jNGSyp6FJaiOsLwQJRjPltIh+PAzUOu7IpDX
sfzaI+HYoocCXCBh+OQJxl+Srs8WFdgUGwO7krKX3Li/vVE7gNJoaO0NE+D17noO
zGdxI1hhHn8LsjTDgTFdpyCd20t7h1rBKbfCBrMcjrp5wkKivZHEOXj6XCgslwc2
L6tNU5DpEEAXxD81ikyhjSNyUrILi6NF8C/lcFsMAQYH88qBKPt/XGWScJdtfan3
SoziSse568zqWAwfDvFowZqFABNaTY5RD/8b89jSKnPVRp1A1fyMgv+Hy/9fX8lz
yzNcxJPifMH7DWTlmveaZ43ZDhanis/Sd/7uxKygsJZK2ailZelAi0BPwGNdLX5R
ioJ4+34TpBQba5blhflhntcshuZcdkLUGhGlk0AFSNkgGWu0uw5l9xpMgQwEcpym
TTS1CvB58RviP0vMG0+BcBN1hiu6hekl/NGweWEJMZNeZOyw56qdYY27Ro96wxk9
ri5W5jfKQNqkjsPoHBL/4Xn/0+xQju/ABjk1pWRkD6oso8f7FzoH5pCZnCGYvM58
uxbT2iS+53HSdTiimPJeKv4wxm6EwEckiHCm/nArG6zNewWdA8H/voOiy9c9bd8C
7cm5zNH8Qwd4Q3y1f7i/ykWy97PmPUYAdBbAnGEbWs9gdRYaDjjlIDhbrQCmwdoL
Poucn0XdbLoGAOvHsSprrS1vce/iok/AmHKT1nm3VDwMbbg8GvH9/42gwDWV9DXC
bDz83aToBPjLCFox5boYygbsBK7Tgl1ptyh/dalQoZxXLvjO+UVpDetxdv2xlQDy
SImgKL+0cY+/kgjbCzm/HxeyRGILHODLJXob8Fm/1+5Mf9+Wq3D9aRFG6S5/PAsC
u1f4LYuYhSyfg19+41uNnTNq+R8/7YrsmXuWH3SOUTVUEbaBDqA8mLDdRQXaA4qU
Msr7bmEc1NFHRAbvb3WqgYQjwCyYqGGj1YkibMyNoN/zP5FR7WpwpdG5rqXyw0is
3rRq03YMHtIbXlwMRBaIhEUZIJxguwrB2Oaof/pMfXqDekxqKOz0j8arh1uLvEKR
RlpUNoKbftfo0As2OiXGbfYSS5IXgJU79p9XGZp+0LsW0wFkU/E3TO2apHAg823g
roLbA6I5mzWmgy4l5JYYyGRVSIOYXnsQFyrat9EOOHxwWoxqH7YHwC3SGOThYgiO
a9+SL2oFm3JY9/v9iM6tqUov0dw+A8Vo43aWD9hAMfT7nN7HqNYzRywPvyFIfo0j
V1dah88ZHDHyeqO1+Q2KMmLhl2t7r45rd9ZhJZNRYfJlr8x3UQpIbVX/g+gceBgb
yHfVZ2pPkESJ6rm1rP4DfXGgPk6CTB16CExBN8vChfQrqPsMtJLUAGULNDm4pi7B
Xr35feQXhjgCgME62vJ9FAf0c3qnD0vXnE4MGwBEzxZZdexTiXcJpYgYuuJPTfss
stSrweA9/7QhdDes0ilRheUMzNjnuEAySvEsCraX5SYRdJREoCdfmiXSrUryQL9B
9RT8WtcbxzeqwJ1zSNBVPjMqjScjHVRflpne3wjdGQn11HoyNcwebvSjhcrUCILG
cFFJIWw5hFRLwU82HbrBA++rUivwstEA7lGgsOWFXWuQZi0zfofk2ag3FlSDwrrI
jjRo75p3M/QwGCVjQ/QqiHbKp1zkXCoTRzxCg5gBbePCV00ZfCyVESrel1y7Ung7
SG0yyQ5OySTY86G39usnrJ1KSwdRjgyrRJy/irBpvZ5fc+z4AHSVoAolM1YA656o
b30M0RkT3Y0UkodGIJ4lOW8WePLtpb7QNB0BBYGSthQd58NnNWkVY44RXWqMS5Fx
tdS5APd7FnLSBnUzauasM4uNVNWmYUkDE1FGHDvX4v79itpfm8wO1pXmHXz01tHw
/KxT/ZBAr+e8gmXCxGEvHJw+Z4cn0dCv1O9xXqzD4ppU20DACNAhUuhZqLMy/DjI
VO0s1v/98JnlCvA8DXVofN2YEtdjey0HAPm/qn0+pOvF+j4taDnQcociGWgB1ENO
FVpc9qbFzpxPdKtoclWaUbEhFXhQccBE+1GM7ULPbZrrM9Ver5gTNvOeUi1odpi6
QnJBkjLxa1Q2HuX54gDNBApXB+ckg9sRJx8k5FZA+pbRaxZ2vxlDWVOBbvhKUqfF
18Pkmyze/gVRGBWANWBXNzcJfehCMVMnQyB8WXjNREme1WjfDoU6gEcbop2MkUGF
mO2pu1guPnqqtbi4V6w+iZtSQnZC2fOoAeSHvBnWaOcipnQuCEfLlCuP0B6+yoEy
/in2j1oe+EZ5yQLV/aabIMQpIus7RUIGViaJc3TaCuWKdGfO7EWsEwpHrJcX5ykW
sF2XfKBS92bsvm323QlKRX0/KeFiGlHc3C120m/K5bghYltdPNCbnmGNIOst32TT
p2jwu4sleyOkFO8HAED+c7ojqnaZ4fUJ54r3n2Bl44yzgSZRDOVg5bhYBTSrn5b2
Q2aykuyRCg0I5komSDSy6FLsZBDbdP6hQwz6jHPYtAJih1CeXbcU7jLV/YOJxEho
iuovtOPSEv8bHowkKsrmMdK1beG64ibz8uTDCPbfP37bpLQBOujUzp93RiDDEfrg
mlIitKTd3JgH7lbmM9zNrDp8Pkn0/XcXOQuvH6SdgAcTmbFkQmRLD8hxii7CFXkG
VIrr8bwJDJk1FHDqL1wAMrkgkFzG8pN58yz254gFQGmOWvO45XmLDSzJ2twEhP8t
8MxuF+udo4B/4pOpu6smw4jGSmTSQZ90pU1LJl6fC8SFKwBvW4sgvY7RaoTMmbTR
xoVT5JRnYWT3EOhfitL2QKYqfsXpNuLshesIPL9k+h9+xiCc1QCoaclhpfaDBI9k
OBkw9WedI6DuZ0L1y9LC+QJ+8XGqTxBNpCz8HycfXYIo6EJ9/AqlMITIXc5hW9sz
Jb38C7bpV3Oi4lE68ZrkCxFwFSooknduu0Q2VpMQM+zgtvNs81Zk5QJ117nxK84T
H6RsW6VP3yb/nNfp5cE5EhFip5aONKvO9Vg2OYi3O6rP0V2LHKd0SCvTBt5HGhpb
vFW/RKfmN6gJrM2Y3nvXvITvUupeaU9q6EQD8pQckziOJ8NUDPc+VS3zfpXWfjJ8
uy3ZIVbFhKsQ7BuNDb6/soJPSuoymvwn1Kdkr127hZyZet5Ky3jgkai2W08/5JSi
lYXuMnApayGmMvbBOCR5pfOo2lQpwAbgi72zixJ2a5JteCD2Cs7usT3cPoTorSIQ
cocv6cUgDai/KJz5zQq1uUVQJA7xFM0lKcHuwA5eSFSKrK+VS8P/f3qfs3oHeR/B
3WR8XEOhedPSuVaRxmdscSKVjs3JLcoaxHgx9PV+mhLaUYPxO2M8UPX5X98Uvs8i
nzvDbsjheTlxdhEjc9m8rOmwgSX/8UclnCAEmzCwPPvLL4UUY/GKTfiSYGENsNCH
U+2sJJKg1ydkdeiqgda/T0mLXefi3zqdnlHh7XUBCxjSXbLXQFh8iLrL1ZFAcfUV
+yyTFz+9q1KC810Rvlyd9PqsUU45ANknkZexdcDN79TXi1cfcW3xHM3cQX5244oa
t2IyWLA4QG5jnDw1oQskYKs/dM9jpUPvYEOpgRFXz1iwnKKpEal1+PQGQmQlVPVk
vM1y/8txmtsuaexVcirFBha5j5z/LaBQvotnkVxEqk5mNU9UA3aGyxxCUdvWzCPX
1fXY5Tg58/L97+xg9HJOaEo1S9nm/jLJcgZhbgCHJd5le/mtkbYur6HjlAqiwODG
zr+Wbgt/eq/hdUmGH7mtXGya8STyFTMDt5xwBFPwsQiTap5YQ6qzvV5CwowtUK/l
OnTYNWj0zth7DuBIHRcQ1ykDwe7GHXl8xZEz0HRL7FJ8g2iSr+BtHI1TFn2/23B9
lJA/T0j/McocxOMxpEoX13/QyTOQVkRFI9aDNd0w8jt31G5yuN4Xq96q5HhpUggi
kwsCqxVOKiIV6+uhltG7TJc5nUHybySqeOwXSfTqtUpQz3r0XHvMxB70tjYKqt+i
f+bf7Oae/3fa3bx5ckhfWcnofPrLrReAvTEKYQYhc0GvVSNUJ7EQcwcI1htTxLaY
Kqog6owzWVoidNvzpJgCTFT/Qyya6Vuu+4qbZqvhCJikuwHRc2Pnxy9rxjzCVoUj
EkxXjq3INqhQdaz/6DFeit3ztld4OIcEVQZMYM4E8wUM0k3qma193GUPm+Q8BkXE
xZ9qs9wT7rZWywmOt5XO6CM11FBTfFeiQje8rQi0czNklt2g/FnmR0qcvzzn5OIQ
ALNVGgL7z/0TR1b5dOnRKSpunYkS/A30ITnn13s0pFFJnls/9Jr4hC6mOx1k5lZn
4xiC9MGylV0oJIsxslAy3L4aZUK+ycIWnG117J5DaIOhZ6/RAqvLB2zqjmDtPfjf
AgwWq48hku3kJT1/EE0WZmqWrxnhvq6hoFTJ47ptQi7PnkfHbjskiygEpJEDSrQq
5MYlvbZQJrcPwsIolGY3cGYHKdyMVqdwrVfqt261OK79pDNoijSDUwkY29GLj1wC
VdxpeaCFUPpMXkYsuAgjVmhVLT/s75l3J80u0+29FSrwhRpbJqDV53n4J52WyfJE
5shwdPINNi3q0jl2YEbQXRhFDJN6gkQwNfI9xUt+fhmdedV2Tc2rCQpb5RgogpoT
ySeyuvcl3lZu2tHX7frgAG56k8lkU1P/fvLhrc5Rozc4a3zsn425GpKkCTf1tIUB
26dlWTeYlSLyasDvGsYEZoFEIFi5kIZPXI9K4EJC+F2U8Y+j1gNFwVq7DW4Y2pyk
xpO2dzIyTf1Okv67sLcveO6efSzQNaIlWdr5pkezAnPkNVoM3I0c2w7sY2xJCBQY
c1N37UbRDfMpve8qiXQLbXH4zPEgWQAnq7A7N6bua6cK4zKquCx7lTL4Yl7DYs28
+TdslE6akqFxcM3U4f8msbJtdlQEKRNylWFWohBWNdTcXSJMz4yyfIRGuyTaBjj9
9IWKP/CK36/DH8rNuwNPcxpZYuASqTVlF+p7lYdJQl7tM7GiXRw1HpCp+SoSSOK8
1skL6zj/cQUYrqEGKAa6IqT+qpkQKuFhfuvCgGtE3rza3ZknA4u1tOapjvd55rhp
0AFGLj4NrJ589oTOgwmdmX0eDUAIC+UKzenTvuEU+9J8iS2kjY6eMhGSv8574Gy2
1Jh6CoAXjH93EaAT3n6ovIKkaThEerqvwa5eeeLWCWlf9WfHCsaniXkSct3sYNiu
P9TdvyNITR4P4ZgFxqAoW5rJSfPAYQWAGiQUB7/4ddIv+d957k0BXqoh8nQ6bwpf
TrmAJ0MmTfQd1DyPCBggt+4N0UsPjfV+ES806z/DW71zIE3/a7jpid7L/nkQJgre
DA4rXaZmtODgEbTnFMDPcohtFHn0w8DDwMFiTIhu3Ec59ImOvZtZNQqiCOJl779q
DGhfW/Y57WoHD7GCJVN5Pe3wm/L6pmTQocNqnmvV9DdHZk9JW3V4K3MjvKCVK9WR
gwcIjbiuzbgA96O4M80Nq2rikgYSouOOxuqkv6jno6m7hTNYDTomf7rdQkQS3HBA
vvF39vG4gu99m9CuwvDxqK29U9KiXsFS9LrxJveX4JlhXGP1oDYY7cJN8E9TBFly
lp4wo9v89x6RQVmj7BPoQfwfTBnyvNjM8uXsfsU/aSH0jKT6mmlogqbT3mXoxorv
cbgwtPyskSzMhv/94Y68gvz7SWPjubFkGjSmHzFYJg6dZvxF+NDLzqc9Rx5vEbCX
5e4sEv93j9yuTPMziZtcAJVemlUgKMJp2JRxPJ/LY9BfpWmcwCFnYC07ALSxxZJd
gdBJDnmaThag+gtawFu+ZgnvIMadxNJLJj7WKIm+IPMDsfUTdAZtkSf8cwpW+yWr
46uxjFeieZTX8uKaf6UL859ErIUkNNM1SDDB2dfaVGKrPPrITXiOw6gOzHCldBds
sDjOhTkVQKLY/ijQbEtGT+CysvUh0xXPgtsiKQ55AMQ60r+5mOMrluvmpbnp9WMg
yXD+OZTTHAOS7B55or0BBOnr5X6O8Ln3k2NqUI4+Fh5ljTzmkqHciLgCKkqDOK7V
3kf61trEBD79Zc9GiEGpLxTJue5yZTCKmdOm5ewfnx0y5cY/IfKUP7CIWnskfKir
FWzBMd8nN1Z1FEAvBVNe2xwom34JgE0NJH+tEY2yaCrHF3NbrxPawRnw5vCM1Vi4
5/A6PcxTnTaxzAp+RgDAq+LLabtR3x/LpPBoIThr+olKhibZRN9RvCu+jkpYYpmf
YJ5prtoWgmoO/nbZQz2CTybyTdaUrHjRHxADWXS/9n6LbM5w3d8J5F4AHg7sVry4
tGNRYLe3cqF3YobJ68e09ixX/w+rBVjm5HGjiEEmB8v785lsX/0v8CyFVvY3nD3+
W3oZxv5AUMeU6YQGpe0tAUBNx3oRYZMDK/+0ko+Ho4ytbnNeNmIoHGKyS6J1sv+N
5s8Sds/JelrYaJ4VLOALvN07nNeKIolQYKd4jtPNGf0iiiYIKn8gZN9C7ugB2Srb
Ffhw5w5zfFeoukA7g/kqt/opWQtqJSCbTjTDhCVpzz4d5EMisw+o9Rx6Q44Bh/BU
1o5CG9iHVaypwhVEmob88x0iTz2xowqz7vxAa9D8qn4iFKvH/hQCuH8axEsBFu/x
jg0bfq6yXrTlcIV5OHRP13K3iSMVyG20CC4kK06PVUDPPWQStOZgy3dkJWtk/PsS
FdaRBS2QLyBZ45ZiJYkRu+Yna+7ObV58hYj85Hx1HWQadhRNBXzs5uYtcPxxK/+6
DTkF4XXJEPm4fx9Jj/i6VKgPtJl1k8WNOYYH4wMa3fhqUD2yvYCpXW7+lK1QODCB
hFAuxjTfe9jBojB5QRGhpuEBt+ZX7S1icukVLa8xk/a7HUOQhMDw8qa7U7iFO4KH
VRav1jOXWVzn5jS7y/0TVW7vpOL5u4eIYYr2t63fQuaf0bvETF6/Z/R0D6B939Mw
wAYyJEMjJf7oNLdPbake8MDB7flplIJLbDxmhJLp1/XM5/QXCGV2gCSyGoglHmZk
eXJfLigF/pYeREvM7OCViIkwmLY6yWRntGDkrFkAmzkRs5VvumBWeef8uXGIvzLJ
dJ4FpNlEfhVKjqZzOXRnFcRO97S28Besmei85tP3Cv+W8H+F1T9HjGv0b1fPAscI
FbK/ZxpKYmQIJQMyJe5o1X1dmCgReB8qLCcG6U6wSlkeuVRcuGdWrTcgbBOlIIix
7Bpxb+kdVhLNIIPFlVXPJHkjGqkbt4hQNdINGxRsd3+0Hhrpz1HmcWR44UkdAtpG
d8m7rOtaJpsBsUXcazODDhZZIIpO/URQaH84McI3IXLLkOeRWTBpxi++EXNB+/qV
xbNFP3G1oPBF6RNdcrhQ8HnWEIg8dP9iewNT1DKTX6WcPorTOS23VySKdYGnZMGX
37HVT96lt9fKwF7n4uDtq6NJN+yDCbH8hB0boBjRo9vLOvXNTQDSzP35O3SJpbk4
D8pAJCrpw0WXq4Gf3lcsz5gyuDN5o/iZQEIkzLTfgfUVYAmULV+dRSk5cBeFdcNh
epj+sZPW6wisWqjKgzS/tdpZB4yh7bEjc6VdPs9DZriACacTLXwnHETXdwcCafGr
IuXeBNPwXEz1fb+46KUFgKa/iRdN43JKYpGYGMy/YN1IPLywDmX0G74X5uvL4VDi
DhcWSyS9vwQNC4zPj7BTTFSNGAwJ2xBeq7WT3DI79ud0CeJynEePf37Jo9L6peN5
Xgs6Oik59EE1iypxVzCIFqxKlMMVLkfy6Szgxsdfz+CDOGK/qqybhB27bdLaS7GG
uz7fXl/J4jkoYz1DJXAEFYOtDahGlahRLEmDLFgenXiA/NhV6DlNGH66YjwUa9Xf
V4H6UElJ6aoZBXClbRTjT6gQapcqHMe5ab7shPDxQRoJIS186jOaMLq0UILvJGWR
0IdOvOvmsEPl4JKogJuxPkEVVHozmrxz7PISDwSPpIitrfuBgRjY3Tu1UryDDvql
Gs52un7zE7FsQkeobrboRWnHWV5c2h/LbOdiHh8+DLU+J+JIKSbznvFpaXhiqPrs
FMI+k5fNPva5F3tBIakzmvAgqSRxN1cwCGFEEFXSjLPvhfWPaYbWfjMx7gJKBR7e
T0Diatwt+P3O3OCiMowlvwyUv2QzM7PgDn3fP89+oRcXJz2ExyhqqzY82Ibti00L
imD4Ad8o/ehz7XA8D/X8plzSiM71IauTD9K51tzQYS+qT+yCpBwdvhFsMfwRZkul
HY1kXpYwHKQHDYUvS3lK/A==
`protect end_protected
