`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
fPxlhNvsE5r+jWGMBCLFLu3yDzmeFDa1cY82HlqX0UeH+ksrMEf+xoqwtDPjv2Kb
wjPiXFJq9ky24+vpEHKgMKyAbybBw7JKWL/NQFA7cV18LzysuIDJDtsK0xeKbgDM
zTLQWyI/I/lucsEaFhzIK1P1l9l2dGZkVoJ35CCmxv8ZZduWZc9FcEzO8zjPswJD
d3Y3wtIN6/IZaeQ1hgptr2/Yvp6jGEbwlRaahBmFn+9fbgfsnKwWGTJ2KBvfc+Vj
FNN3lVBDd5xGl6qmg0gI11Tukp2YpDHe+AXPfkShe0kDtl6pp0uVVxJ5JoC9eVmM
xLIzP44VG/P2xf+pbWmYlQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
XLqv1rYFC9v8/8QczUf0bVEAmHBbKnMV5TTmW5cfzAiY92/EBhBA477jAE9aFAzW
BJrv70EemmVWrEG5QBJ9VPYGl4j2Y3YCCVTZDfXL2ePJWU66hhLo0/QKha2E673W
l2HoEON8qb9URZepE85IEw9GkqV7kEMRs9XDknei7aQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 39840 )
`protect data_block
Du00/SFz4JWv+zYBRbcoQf6+cTISmrVEaNILAILmDMz1S3rvf3pgAodsz3gTiGpj
oPx/NsRtL2YogWb0bM6GiLs0y903W23lGZL0Y/wxcvZYc2W+gL4slQpRLC4zJiXC
PsZqiJbkYwOSLrv0sDnuuO0QyXpKLDT9fFDgHToqNXlxdjsI7JvxjQIVDYI5AASi
TQvQNKkTLl3jwqw5aXIutlwpInOlVm+dIhMkdI8eSDxmw1d6p2lSw+PRtf3eTzzk
8meoHDuusBLfKLQVjCdtLcLUYpOxD7GGAbu0gnmzJdYnWLQ4CJXb4iORASD7zQcV
y7yomR2N9IJVB+UvjX/VwEqigpQxPEkChcm6NdwJuUuNHGZDEo/p00O5VjsdKbYD
L0FCnaaf0uv95aoLxmm/HEedd5HehBYSaepBQNqTd0WArCIVrO5S6NtA0BcMBlGF
ymwpDezkpanuhkAhgmpDcIqDtJjKM6kpppNnbQgpltOoD95cT0vPfJL98ZGrFWH/
qTBPaC5Isio2OSXEu0W2mrMOvv/pN/ZjnhzxpDjhjciX+WjjCHQ5YFCpIyej31HW
KDhVpFZ+VvaGFM24eioLa7d3b90SM4iL5rvm86jmeoZ63Y7m7Ym9EeaoAN9ih1j/
fIS6IBWwl28bIyUMIqJQI7uy0JsFP11D2yVz3MxCrputVJTW3ASYkU99unD5x8sk
KNatH0wSIp/2qhKFU1VyguRmkc56hEtLHxRqB8msJgfwcsLVnP95BRdDzDS3Ez3x
ST+MUEYeklWO3jEufzTr3w/yBF7Ce+y4aJerh5I7hTKnQUfCDMXhmunRp72UANuD
DYw3xZv/LOfPw5QZzyBnVMgRPn+u4kbWsvu6JlF730cA0Pm35BMQyZpEXUMe1jem
rsVUtkTjY6T4LGLKk3xYtcAOBEpEjSObt/X4XddjFftDTpiRGvFA+XpbdoZzSfb0
mi0tzj/OxAcE3BwoSTWyw5p5rjAk8iKWEbYH7UnOdwYmHChUKvhaXcldVtKIzDoa
0SyGRU9UMbZsE7hYJA8k32Obs31CyRUou+ain3wY+FWL2j8nRXR8J7kNBDwo+7zR
pgC/ryD1GlQpqbTlOzu7cGHszNEA2yVA3UP4N9uTkG8bGIpA40pcAYVU6aPYRkHy
j3Ks5wygU+iw92jxY58gfRoUSsO/jQsu0uXHKkxs9i8iSYVlxJZ/ys1cYJ3K9yYf
YgTnl8/l7RQk3sV/h8nhOLjzxZAZl2q6sW+56MfOy6Dh/XAflncIPBpElzI6qu/M
+nT4+c77C12rCJCqW6wFNLKEirz78Q3TtA3V55OywjDT93kLt223J9STaW4pDQsc
rbLJg4uN0BS1e7WkLN21sLMICWFjeZk7Yc1B8S4LcvuWuifOJRiWPMdHzIV4Budw
RcLF2PWjQyoGqJbT0ZpOUSDCcq1mivCqv2dq/f08VhPkC7vAja/kzBfbK4rICMii
VcVVSmXY5NtGZ9GKzfCX3otnXx7xV7TofdZLL9iijoeMUevawc0a65QM/OjlGvPJ
9sKumhhVUxkMjiK+RAvcm8c7/ND97bw+i7PrI9KI6Nf0y2vBmP52XYVv2+DMdS9r
SkZXAqmnNgv9sRloVaTKq14Q1HqDpIrjcOggwskSdKT8RbKp1hwPpR3HPoQKEog0
dhLJaJcUMiQO7zqfEPX9g6v+CKaOTi8CovKANAimOE1iThbiLM9GeHXo0fSN43Rl
wBpX0Io61Veiq3vLh7Kfp4d7gdwgxrKWfe0QpPVp3a2slKZMnneOxrd2L1/HhxSU
UTY7ljl8BdA2ZalVh/nHq7yIjERJ8uT8dmOLCEGFarJnT55vIeZQQ+ImESJAlRFX
gx5FafN13uFjTHh0d6LysU0vmXcRx56KNpdeaC/atfq2mBDECN/9kV7hPeZFFNxd
JJZmxMG7d2iOCXJs3wMRDiOUiZJh0c3urqtJsQV9Mn1pRsosAidDYWI9qsYtYuAn
oShPh/+MQFwxfb7NaSvVX1WdOxoY5iBkhCJc0F0MTPUdZa6Pjpc9Q87qlf+408o/
1BOafVRTC4T0oYreL8SXcVDMIey6WfVZ//NaO49rwEJZSChfBS2fNs7hKWLiNkQf
DaeBwb2NHIio1JOpCDO8lL/I6C3Lrjvru4Ky0LpnTflKa9jqbznaShkIoiAehvI6
4oqpI7pshDiAj2p7d9jgrBWcogyw5zCJ2Rx6ky0Oxew7FeopfeO2A0nZi7NxcASU
bOzQCqe0t3KEXpUE6rS+Mwgu+AmRC+s4J2IzTzmRiJgC0Au0DGDga2QnB2P3WNHS
RbWeQiu32WC6ifDiMTmQmZs2wlj+DIItKakfj7mhHw4QOOYPp51GHhrp3aUOxCRZ
AGRWTO3W9Xyvwka4+O0ouq39zRMcUT32m9ywaV7nHRXTjLrAcdFYEi5alQxaMHJn
9Zg1v4JFQDZMQ8fowdUmpJ0ZMe1+9IFJqySx7pBR5abH6f/Ng7YBPVtxNeppkkII
9Ba0uGlKg05yz2jI/7gDUtFxpHowvoKsLPjhQqtK6gtbxSEPa6Ix55ttHh16GOeV
2Xtcdm1JUG+P/0kE6ZcwfvLRSbUYNOSi733xV2pGxwhftc+ix+mHerKFXbd8KqaE
EvJV7fq3bE97iaTy3/5v5CsaPzXY2lAEHC59Rl0crmWa+Fv6+q1wCb01uMaIv/h+
mQOMOkkY+c46qdGVzczbXklhuwqkWOc3VcYf1O+M5nhHmLhLo8i+wP1t9PgovPSM
YGgUmY3ciRp9y2x4YSl/fkqcanbbm11GJe/0jckef+ZX3WONXXH7LhGhT9NAoUyC
cFW9idslLwp7IXNWToaMyXjZDKqTfLmYQJA4yEDDtHZHhIWNw+CfrQAweHsN5r6/
v+AGzsAuQzxYrlmW+g5dSpNWlpL1O/GXAccRbIH1SkO8YXPIZfZ3bAGeHRfvCiR9
0bnMVM0vzEKhBaZWdnaMC7etmOUJZsdJN2xOYEJFw57vOxtnxPw2y8V5bzx03ONf
o3L1fDNY1KiJKePMIoD30rHjIiwNj3ClIIdYjoVDn1bJorr7K0qkEmBw7LAXtbCQ
/J6Z+5d+DWlOa8xCmTf7C8KV5LBvsYsKMhMbc4wDp/lIJySl99etncjHV5ks0cuU
uttSGzD+xPSJ/3dVR5xSBkoJWg009isJVcVnu+xhY2TiJFNUQfd02Ylb425czPvb
tDqTS8m00TBgE3tgZ69slWace23+Pnu9bphQcAcvdG9QtPwkOPD7DeGrXB5/utIZ
IAxjpIycQhkuDn+yauNvlczmgd59efn14q48u4fyQAWKY+tJQB+SNzuABpa6jOD+
dNAVvorlN4cBSmG4M+My4EtxIzDvBMhlb5CspQmKidy5CGhbbR3fQhbVek9Zh4ka
Bdq2lq1aSupg4FiC+4nK8hbdPT84lMrG5WryrqK88vFR/ELc6v2RBsGvom6TuokM
6YKYofqTR7uTFAzQ+FtV6VnK8DrTLMEcky+CZmpulDtcbR066XE1yml7wqpqWKPe
qUkwFj/EzYfnAFWHpaxxV5S340lI2dNUz56A/cLV7NS4hTo5ALgu+1AweHsPc77X
emjpcKbiS9lR6rdjQvel8jcEMJVToqTNTthe7UQ5A9AOa9pFuE++kzNm1awzo4xb
Lg3YFo3i2w8QZ0cpoL9G5mr8lv98DxeesxHkRBmjxSPAGUNVfNhM9t7zzCUNeiAN
wC38BwXJ71LcgaP4ppHLG/Qce1sr3ltpBGFsIDjteiFiXPwaB6PJsb5L/lCUaryR
XfwI1dUpyEBtOcn+pgrCClV3woQ7fX5TGyNQeirXjfUUjHXrkNnTSP/EvO5Y+spb
XGZu246GoL+K/LUm9lX2GHV6uAPGLFUDK3AMCmPz1sNyA45/OuRHD7NpzwG9G8fo
hFCgtYBr9OGzweIcJOK9uLQH7tpVb9yE29B2FR4AgdE90nj4cv9GszptOw7OCe+H
P4tMw4+lCyFv0LaACFEhnocxvqyQxLp0CQdFR+95wyjddMJGChKVHbZobUwsGgNf
RAs2268PDtl3lcCeY0xuzgfIv08xnATFb9ZoqKEUJLSglwBVOOYrF4xNn3jOL/nl
tdKpfqMAZvs187QsBoxgCLKqaC4pxzmD9yb1XAW3FdegIllEAq3rvIuqLinhgbxU
rDl2pDgDzq54J8j/WAXrzQPo+VI4LbuFiBWvzU31lRUpeROwHFXJr/wvPSWudBPJ
SzOxIf/YnVbVmklYKLPc8/XMKpmz1z9XZUCukyYQeh5FhuG49MNosC9YLgCd61nw
FdF+S7rkaRli6QF6qUrq403Zr2JFq3Q/vvfiR85Zg5jy4hIG6J3v2+R+Hl5KmHru
5tn2ZBIh7a5oFwHQYSPk8GgVIWQ5+AOISeYM9mYwAsHYGiWGk7Gw83aaQEgQGotq
1S+2wnRekseekXH/zNpbWZAF79dszHKGlVmX5OMlDQSRX9+8k4kmwkjodtCsNI25
WgDrKW2sRKgaDYEVv/YWYMBcJEeGfJY4MDO6a6avWf3SX67ggDjOq7JG7Q2gWokY
gJwwFu9PBGx9cAX8Na5yxqsDnRYswIhSfybzly6lwSauy0OHaoE1rsmWK7YYrzFc
BSAfx8OaW3gBa2jm3ZeCp7H0z9gUgTNBKdYY9ZlyeDEAqntmBUkx+OIpP6Qpq1wH
N3/LshWIys5qKtbiwDMRX1q/mG37PnkpiaFETz/CPO1peTQtw3liAuUmjobB7PlB
B2kqfh+rUBl3szi8u0HcC2XIzqjQ9cHW+BF77Akg2Uoglwc6OJOcgvTZEAsSSFyB
kH5SeclUzNtCjF89JyJXRZWPoAP9tPAdcz1Y9XtGdjPKzIqMTM/pbjnplgnDUN8d
4rAVobueyUw2iXS4dwkk6a0zRjQrn8SZ3E9vz1qHpFf9cIw3swh1o4rsQMxjFQQk
cQuKE2On702YaN+1ReHQ/pkMSbCB1z496pE5XRs7ToXQKMXw+lgYW9LxeF3D7BoM
dXJR7R/omAXIVw0ojigtGkMk0puzAnHh3bKrhHBpC3IIxDiuHAHUXaZGkx0ZiXaq
BLvHKbl2wxEOd20kLn2LtQ8KuKUs459vsthAKmIXDnBaji3tyaHXFApngCOyKP7d
VN3ARe/lwLKpVfAsJyPRk34GdqoDzcDIoBCypYjtR1Rq5bh91wspO61PceVWKYcX
ECGGn/n+2d/xCga1XkO+G0XLIqqrvnPFZS0Iq8X1VQJZxI2MbFEB3CA1a1xIdMyu
pkBaENI28uZbruk/lD97P3u+zXx/rea6z9t10nZ+5vLXmBYvsvLhbvXCC/zs+c8O
zD9OUV18Ol00G8k0uQJq67LI0JPKz64KoNulX+Ir/Do9eSHwnng63LMhgUKdB7MW
o0SQ7lnsShLzvm1N02rpiDfnKuzSbCXaJrKREyOrKDi+TA4N6JQOss5h0Duiml9+
YjI89MaO2Z+dc57BRWFB+BsMWEXdor414Vo6ydnfPMB9tmohSU3yCo9i+GDuM/j+
2rP4H4x+OMKldCc4JbeVBROtlMIBLRxUqJsI9XRzUEj5tmzJgWVe+gbTU1vlBJWn
Xiht7kOVqgYaCE7usAaean7QfrAIHbt9GH9i1buQPZAoRpMSKwdA3IA1d9VrKQmo
hTOjr3XgpLLzp0AvzDArvJQnM3RF56vL7p/wJzsbiwBo9LrbXOFO5Pr2mZsa90qF
bjwf8TRS11vfJLSLecoL3BlAmz0tbdg8dh5fJAjPVSXvj5/nBwVFi9s7LZvvsY/r
yyfzz5q0CdaVHrVzaD1FLTNucEVoPdkc0d8RnjQJAIhbKkkHKzPG/IXZnMBwgL4m
NnRH8q0IkSq3LmjsEJe6g9J3Q4QGI8B1zYYt74PEijfKrEU2gA9Fm8l9VVdBIxyd
PNf7RDZkaFYhnKEH9UB15c3swsEC3lkhZ03twZEbX2+fF0jYjYxXVleZiKeYJ6Ig
SM+DEPIko9NqW+Phn4RJpD7IZb8KJQfxkwmHYFM+H9jUFE4dIODj66HOCdvYpHsZ
twpFY8Jhi0W9zfjBOUX8R9sS9xpjP63rDhZKcPCCIuQ7/oXh2Mr5cpeyxdeTPD82
4UwW+2ffiinFDiFIceYE2IMgxRpw4kxsbfRbdJa2JXb8FtTLdHEtX995Ozn3RcVq
YDcV/0R+abhqSTzScN32yr/bsSncp5o62RhFxrZ/PDMnn3h7Hn3b+HUWbbeiKGEI
rI6/amtU9kj0lezxCgxQ5ag5QkSCeoLjRdkJrXcSN7clCXZi2ue6nCDI9GxI5QAT
slJqaQhYlSLN0z/VvPKBhJABb4hwKCIJ11xMJf/AdBRsi/J4j+Kxty5YEDrCYyHJ
r/UvgdyINiM+K172TI80HsYlK2UYZM7H4PgVspE5xapX31J2cTYA0dxEm/JEPNlJ
2pFvLWdledJCvDDYJ0kGaZT53PM7fxjNV39UOhxcc7LrVzn6QDNyUxpR87E/qUGp
2ONfUHJ+/YrTywcoPuwmOK3o6d47c13+4rwiGPUfwgJzRORm6nuR0BoFzhOjprUc
YZEDRCdQfVh09O1JDwxnzEGGp5gAhokf7zSM29m9amT+OL03XDaebeZdaR8KlXvg
ziFiUOTZ+NZanxqI9T5QUzrkuGfKz0L0bXUEKQprJ1y/CT7/pp7iosDg0OOni537
UJoSMVX9UJFNtAXbffvuDSK1f3azS4rfg8VrSGDZBpKcctl3QeSvkWlt7NLVMHzF
8gEtkGLgQgM+qCdahllymOtLEsggLr9Piyny8lS2nwXOajHr5X2GoKMHtqKKkELk
RuQtelTuEfScFft86NBNU+ixpKOooslRUrjIWVka156/oh0irrGBv07qJYt8QfXA
m8Vl4Ey2qA76X1St2rmQ4lvt8nijM8CRxVhzIqd1G9cKCx8NgWhbrqrkRQNWQsZF
nHJU0YdRCvYKmeE/oOnL5ROwYT0kJ/KsoVkd6yFq0xCYMmrsU8mKs8zbOvdSZCKG
XY0WQh41qL6n42p1VuXlp/klPLnWwYK0SNxEbZ+lBSJrbuWti8O+s4hkAh5KEp9x
MTAk3cykHdaYn3fbAS3F8hwo9gFex8xWm3v2db97EX4ynEN6uK/b8ezbZ5LhoNSp
TePL3/EHuNnCnwlDZaP/8ezhIr0LnxMUITUbDUeUw8fqnEfmc0Kt4xlsO40Do14S
kjYbMx7VNMjoG0kMMXHMtMGl82jIxEMD5i0dJqgWpI+G4OSLFqCQh8HhIht5nrMc
1oZ/lKgiwWpvz2hhyLUve6+TvnU1i3Nb8BSfdUM37L4aA55CrbKtxDFwynJUT9CA
2Bi0rRgaURzfOQi5ACV+ACs8CWr6AkZ60RJixTQypno6Ed7pDd3fCLNtooaoFSbe
6HwYxIxdYGbs3czd0oXAy4CFA/pRPO+WWvnRdF5rwtAgkbGx1fS+LMUlNLqtRgNL
RynxxO25DvvOp5hgyLUG6AX4UKd0Uej8OFmT2BRVdaUG23wvBhMgHAgzpZnagHXz
5yhjUc6CeNJPci9L30BwHnhYsoeM3OYzEApDRFwaIRBrnYg+KQ3XuqplMsXfaar6
CPX56aJkh82sN74ru7GPwAiHikpsTQtFoMQpcAFTZ+OcSrKkPSWBwnfHHY9hv9Ac
3MIZh7yWggAXWVv74XcBQ6JpLZA5KYhXkA+wtRaRr0KBTx8I/6RNbtQPD+/aBNHF
6QEFO6baZQVGoT+rv75eXyX3mNTgO7/TuL/A3rnqQmNkBZKNRtRCpXhRAbtbI3ZW
vYRmYwIjq8qbF/SLE9K1y6/uDx9JrVhX1sYgyoqMUnOBahggxF5BfEIl8aHh8vB0
kt2p8Jzg1gq40FQGw/lO56uRxLOdgueazmwWAPEdpD2akKzEgXLlOLs0Za2Pxn+e
3u8CzKnJbt5VA8Fl19crufzQpcfBRHV/miOLojLrHGt7BNlvzszFhUmXritZsrDP
R5psG44JansgOwjlElzBAWlovr9uSufdB9QNdQSSPyEHum6Gv5mEkPpo8A1Baifp
rCH5rOVtjyqm6PRrdYlgxP11ymYFOaMKGACjDemV0ufdGXNeT7NzSg+M24tDm14z
W20twneZm4HIIUJ9rvaexNIOYU/vzgd5CK3N+nCUONg6tv9y7tb/+jeiWmXzsrOK
aP3SPFEb7ufn2tshZ432cMBhiV//xeelSgwJrs8YkaBAhW2YQ6QejONfrmGvNASA
Yj6v3WPokBhxTDAMxFg15TIW6McVmJjtBeU+ApMnziQFQsrrrWWC+XDQrQlpgJRZ
EOD5z7lUt+FTg0Kv5zOdEnGPuJ19K/9lprenVu3hHiiprb+xODj4Mj+x+WTDSD0s
c86R2SB4VawveDJBYicYXZOX9V1VN9BBWNXHI35qy/hm1Hvd41rlemVgBatVxUW+
PPpVcWnwxVj1anGn1OWstL8VDOOZGGMYm5cAzxedL23JauDqi7kZr+9FUPaAyHLc
LCzGNiEscAqe/r1+5nN4JHr0UAoRrj48uIX2jG2FVl+lbDmsEg3kKHtJMD8MNJOE
/KiK9Xig1ZZ8z64h9suy5hO01SU5dvV9ZUGPPjA7VoUxgwQbl971292eS/dq2e7H
GTicCw+SrVpBho222vmQR9ANBeAYjD5aG/iNwvLixJrybiVfsauLbWgza08DWhA9
bBbAqf8ozSwFzs58EX38jctrXwEOHCdHJ7AIHbzH1r4+KqDFvWvv2d32+/JiAcUl
+wokmIMjwMRmB9XIoS3iZ7cpVd3FxP4zT7AXEKNG0BPpQvMCt3s514ENtDrqfGpD
Ep+oc6xUJFjMy5uqvn1MeZ0XXYW/nxZz6+/kWQ3WW9Er1oaquVMvGFFxn2zHifhs
9Yz2Qd55p5xBo2xwF9nc1v46avAe6QJawLPfdWvSWciJHDfUA9VqvEOFWSE7Feim
pUDVJS9X6OTv4CpnrYNgSSIRHax1hm4fPrWIqu6wN409islPjjbStICi/WK/96Ob
w0Hp//QRL0VLMt6/zKtCqz7sH+7SMz0G1LFOrhZskCHYwo3JHtrzrsj0dJvSrVDc
TmcDcKlBhK6rLAHP/shHbbSxNPXcY8frXGd0zSQKqBEId0nK4t/Iv1YWUFulY6RM
IY7gEZVDCVpwXjlGtcUZoxaEjpD5oJQxpt762PbmY4EW6+BFWb1FmsspeAIMBc8X
fRnSW+TO+XyKLAbIp/ANUWiIfq4AMAra0wOCNK0wKrJZhpHQE1sld8mu2C3Kwjlx
URMsuIMiBovidZDXtC/Edqa2zAvVrBLsT8wubbOJoq3wp1wJoWsItPhsosj0JOEd
GJkq8B2fXi78Iz1x4ZQzfoB8ZF5jtSuMS00BjBkBmHPSu13t+aN3vyTWoOlL2VdQ
WzunFsEuAapU/XmnmLxo3Dc3tpSEjIgWiZgCC03wf8jgnuKXXWjiQ3t1QIoQYakg
pp+qlkK0eIe1OAbTBiDFhJNCghpAzCtxXJDYsjOEolxj1o1jwG7TTQ1eGsHJP0N1
hvfSrQeOpPNHUs4Ja4oIYadLcB0hgpIkzmTf95rnNUgHLBrXOAIkTFfG9tqCa2DI
BXZTyM7e6NUgP0G58l6PAX2e+pNi49wXTgSc5QpMF1gXz3SAmPjZf4Obbqo2OMSP
y6LTYB838I3X9uvOYRTcd51P5y2ObDoZnk6w+p/UhCpeBQOeNd8SI4qbix4VL3jt
DEO73UDu7aV+efgJo8RTjBzjZ10gefZpY+Sv7U2TPZIf2Ao3ymfqnFGzNX12cjq6
IVG6zg5Q+r0QGVm51VJYmFrE5Wkwg9K4NKAXSNsMp7ic7KeU0NZyset1SWdjC4Co
o0m0t0qMP9l6es3f94cYS8I3dZirNALxWoBLGUUBuqWnzEX6DfqAymS69U4sEeKa
ze98ILQJY8hmkv4KtBvX0Zi86m/3c2F15247spKE1mwIpz3isrg7OxH9kl9OuftT
ijAQ59FeFEBYnkPJa/m+w71V2BhEh7xBMKzCceg5AQ1avuy60RLWGlNKvdTcdGYO
oDreJwuh8m27iD9aWE+gC8X/iqxBKh88PwFtPVjcCxXQO7sJMP94d0Fa6Cg3bhSD
YdXpyNqYEbjiuY1BFdhOuAbxHTC//hOphOfElLssBrOvyKKP0Zc4YRt+/kiaUtsg
ZRezbkST2Jbt7GHJAaYhGUWGSoEDrj5Clol/kU7h5GjR9vU2dG/Vkk84xmjAt7iy
KrHcO8dgqbuFI5hi8cyH8AjK6ScNIXonMym7tVeBIcQVFxgdlEUMw+K/pp5SCUyf
3tqIyjkb2i8CX8Cl20zg+nQjme3xpw/eDeCHEcRQZM5XJaQFMcpIEalTTyaSSiI+
kyMYJyBj0D+iZy7Z9Cc00oZ2CaMK48e6JzbZxsonT+xeP3bx66UA40d1P41GU8Er
rfDSJ3ZAuVa0QilludpArPmIUwEAiFpRnH8v0aTbLMjsuNxJHRrtEYeCgofPFKpr
Yyshuypgl5grYDORhkP1VoSWrYHy81Z6tuiHnPxpXjQ6KHxX+OnXXkqU1mcZWgSo
LMEBWQkrEYBDm4xKAQg8oeRpfbDJfdGiMi4zKC4xcnkxUEn3lT9tymc8gw3ah32x
DmAxUROXMhMcYUFwsJfhSKz2MEvrS0Q69F+ExcztRTWg/h7g6h4sfXuB1QyszrSw
wApW84vK93HRTxSAXGvZ+g9xnYjQHHV/opdswCY2u/3AyUV8qsB4qWKzfRI+esP/
pbEJauGGk0+GnbFl0b8/qMgrgEZC3kaZTG8BRnsRhCkioFnCi6J2MIdIyAG0YRb8
+j09aBc0Uiabi3BdCZf8v8PrPEG1QIEYAdQQE4jE0oCNMUdBOg/ab2bxLRaX1WJo
CHEFeRbNhfbYf2HQyeyBqtxWzWaqZAl5ba4AFaLgwnSO6WoQRMu7gFeadFSAzMNo
d3IiRS3PAMr6Zs+9+xMhsOu3c2aICPSYqHpI6Etr6z8hOR/FPlQ+BYLR1rNPxo/g
bNEGPvLmAne3PofObbgi/9V3Jt8v0yY3R2gwsPduQR7FExWz3vtJJk2yYk3WyLgP
B//h2n8uYSy/k6fH3/gEd8/kgJ5FQTMRFZQsHbq0fn3f16bRDapodVCItqLFxH1O
8sX/eWecK1InpVf3LDcP9XkjdaDige7vFfHvfaZ6nWripfWi7blWnkRnbvEyf5n+
3H+FnEaOHPNRvmAyg/jabLgQpXs5ilzB4vMWIEQ8S+lKbnPOXmy8bRjNf+89aY/S
mTAGNsAM3pwpM6DSYTz+u0FMPHdmaZhEbZMl+iT23uue+kPBr03RdbYUGPTt3HZc
OG/S1KxTlV0CxtfeKc2tzMDcfdqnyCpugd+p3P/mLOsGCw1bEBBCE1VrcETr5PpC
0Hw6pJOruABaeRnKWn3fnbJKR/83+9Niu3f9XVDg14csselYrzhKZmV8nCXpl3D+
eMCGNO4EKDUvaLQWSfPFWb7BfSo3SFsHXZVx6eg8KLFGDuTN1Us1kuyks3NC0BiW
LCWMsCKGcaZ+T1/fdivvftz5iFKFfNuuIha6R7NloKV6rjJhw5sD3pkmKIumhkG3
oFnttqWK0o/ndOqnvZnVK9/AH/wyGBO9zDDlWuvFCYn/EBuOhifRPgYAXPgE85uX
zZtjgH1P+ccgVEezYEm5Ph+9Uh3NbmL0E3+oqp0h2IbYIOmpBZiLdsA4z8ZcJ3oa
DMMpMfQW2NQma6eh+K3n3cRKq6Mdlx14P2brOcePZpnrssOe4CffkNgdn0wcSqOj
CRDqRjCbMsB2WIye0wNVEDiHhczmrAHHxormDKVYV+uNy/pU2dsIf0hFjbIngQIU
7nkkOgaOvzmypcY+uV5ZxEqN4HDwBrnn3yiUBf+P0EtCiWNAISerJ9F9jG9HTplr
Ynjx78lPguX5EWoNm5gJsgh0QlrWA+84tonVLX6vraY/APs6S0GwK+Ok5kbS25dG
Fa16jUKBxizeVjuIvwe6k4avI1PLmeF0S86hQtxduLzLKhqYeEW3lMpJj8HhVW8U
F/Bi0OrJXU9RlX+A4ink61XMk+swtjjCXrRrO/oZGJtpA5UgL/Cq8v+fpCYA1Max
xfV+H5ThZPBMwYAMXZoL5aEKoz+zp69Q7u30yO3KIt4LwJemZ6c2o/A1iNZ76hd2
QT5mL222pp7bpnGAueQvJg6/g7Qh/6KAbs2y2Owbpst22fcm4QtGUgkINwYL5oUc
wHAXF3LIm9ud/MqHWyZGk1CDeQRSbNpEHr3fDDP9u6fCuS1DqD3V2yPmCiGx8J6V
UelkZRuiSTB01XdJbnY+4bq4A0sluGZDZjhzNdQf8/ustI2MqYgRFFUN2fIbfBnV
uuhwzsVVX56NIE42ZAdU7TV/Qf1/7VjLy7egKyNNQ/iIkDvLKfaNgmcNkGJhMq9m
K0QkCgfRLDDF2pdrSMHdcrDcs8gIGp3OpnNQik7ae7YDsId+sp+4LkYGhLiSjtyN
eLNQG7oXPeWzXGXqyfwUdgDbkpgy0fiSnvl1QOLzgck6vCSk2yzPUc22SH8kpeQS
mTtH/w+/UnjRUU64U5TRkFlA2fw+BREAdkA/9PMgxeZYSC6Z6cMdOjLFb6JTSBDm
UoI4ri1ARfmF+++YNdsho3T8IEDWehN4M6vZiginU8BHc861BI/wGveTS2NJ8jEC
1pXDXnaQK6TGUyOcklpd1K5GhaKmqRVIGRsyiYZIS5GFhNJ+rAr6rKHNjaRp2Q2k
YBZ5q0SnHcjAL+y/hwHJ1EudLwi2a0LSRxf+qqvx7ugY+yY2Jr40+SiWS+t1st3w
y+bDg3y72Ck23YMeKqo3T4r21EykfPI80WL57tx9RUXdKx031hKqDKsl1hzRBUzp
uSGdXK5cxJq9/m7TFx/mpl7xuwgo12JM2axRUj287xh8WTw0ZPwgOQJ+6QZ/hVLR
TggMbIB027fMkbwaKRvCTAvJEXjnyzc456Di/7CoLkF5hVZGPWgIz7vBbL2qJESf
wkC/pnhvZ9001jLIU7cxiSZ93XxhunbI4z9csqoRypFodF4UBLuKlNn0RaTxGF4H
nmM3bgwCsPuTXFabrl1KbC6KQxJl8AUi5mE3J6ofXagPCCP1LoLxdb3oxDK3YeyQ
fpYx8rDvj2RoEpY5yec+IKO/FRk8MR+1Epauf1k7nF2qSg+esCUrPfbEvTfVE+qO
brBDCDkFzIMQU4iVR/qKSUwDy819oikSaWGb9pAx8bOX16YIHHlC9Vu6BETBSIfS
Py/+KaRRHwNMqm/iDKKRigCa0emTZdXeslojEk9KCB63/NIDuG4Vp0LVdiG+Uiza
U44C5rtmLfkR6dBY003EClykBPvOckMrDDQl3PkA8H/WWMfBZwAxN9dcaiglfdFn
6AM/vxr51dRiIXfPG7bBdxIiRVsYSHvR4i3TNaLfPgK+XGJKeWigKrW5elUADG7p
HXys8E5nIvCACjmRmSoXx/KAueiSugHVZiHAgU8eKhRE+9/9StP5HYtjvDBahM/W
J5+sKY3YAYE/y6g/fWhqBm+TXrG6DncJDcR1LRVB23zb9PT8k/5zUeDRP3n7f8gZ
u8vj7WJ4xbyC76VwIWJnb6i+bIXdnf7puf9hFHGjLFQh3SgUbAewgGC1wsbQVobM
rDQ05+vIK56sNonSNmhbg+f/bnspmIW+341iynzjo0XuDAb5EDlIwxZOyfDOcbHj
+BjFuc3QgYBBgN5W0yxyHpkOwjJ4ySCfs8wdzWuJTCTabolr5O1eOvnPJ+M9ILFs
ffuQn0+VGLysvz7iA7diTiyJ+/Ts/unQ/Dq+x/eDII+8KL0aJaV6Y+As1jes7bvR
lKHFDudyuF070mcktLSG5W0QQy2ufWc1Ws6kA8uvteTD3OBNG0zY/KreI5T8F9M3
bYW8w3tgPeEN/PDnnpcdhaoJdxCSrUCea+57qaZmOFaCaejrFFLfX+37JGyIv+R5
Lcpy1Jam5idr6bXEDP6nF+l9fu0zom/iLNsNNs0EzKKWvIURGuJW6EeLNRC7eI6m
/xt4p3niStpbkGlvg11M2FZpfMTBTi1kbcDOqa+Lk9NixINeRH9V5GZvLMJjMyVa
rzf56Svyitcc/egXOHrEgMMHqx8Q79kH8TJppV7/g+hOBky/PABMUrMCZe5BGdlc
PdkYl+iCJBPlzt5Y05Fj710AH93cJxxjccRcRM2Zc3xgJUj+vnVY2vZ9lVMWPTxL
S4AOgDWk7+uBEWvZot66cnwXwvxYjmbrZa+szytKwoWkeSEW19sMndVKtWFueHsF
dO3O/686Ned+TvPGQL6m2aBXLX4zlAX0A+Xae9rXqrEaWLaXF7ynmmxXPUyG/4NH
ah7mbo763dssV1/P6RWEo8jBQCDI+ZjgVqZTfkD1epRrp/D0w87JwAw9TJcfjQai
XlxofV82R3Ky4GuO4RlXz2Q8Xb0g5vrPZkVAPwfeIA4bFm6pfvqEHeThZKMNEi0P
VOtLFToQ+XBmNWTseacrUBKCdDpF8+rTS/zTLpm+wFtb3GmZvL5KO5cutnaCTmDg
pYpBVk+pINEC+k86Q0dYVPq9zM4gkuIpMz2sNQVjTyRSCPSeD3zvjsumVp31zfH/
iC9xvq2c242S3Mz1WVz99Bk892v9Wt5qSB1Tyc+3boq+RTrC9dcBosehWYYCpCMS
lmxnral2LSD7t8re8enAO/RCOevMIuxpBzIoiQkhQzlsW3XRkSKu1ZQzvxHsEm6u
Gei6GKMX599KXaeAKCx6q48RxOHcyNvYqXwIIE9yE80dcm2fDq84ycb/baj0DN+S
FUhdu6biiqjc3g4ZTEnALn++AtWFp75kXkoVw64xT30kgPl9lfrS9OfCybKiMTyV
qJCb3KwC4nLquTVmrpiDFgSjMM3QE3zyfat1HOdazR8zT0Wyy8hDGf+B57ehHGjg
zvn4/gfdh0TOmwGigBi5jEH3L/c+WwCJ9FftbGoguBTsWGMhza0Gdvpebp1nyjpt
m1v1X6IZYOd/E43aQKuu8MJQB35P8KXQRcH0y0vKj6kzSX4STkYrna+WAGz6iq9R
cB8O05e9+tEiFtzDlS5aHROEGIsibtsrQhDrFqEEmrJ6ZFLMpS1SKRadPnX2IWkN
J9I6z7TrdI7H8hPoQoSziA0PForzcJGXcGVcdXTXI6U+edKcvAcbuROOErqXShcQ
UxgXgGWeGKe06C3xSVkVHd8HopYf+wvxa6vZssQZK64xEH1n/fl1ewthLxNSsPOK
wfEAKJeY0UtSw+/ja3jN4DCmZD4EUMtdjQ95cArR1M9jcvCU7Qly6IexoP+O4hHH
iItllmCyFeqCXgncp/rZvqmAC+1JBIQIc6Tx3Dp1nknHDvjqzKK7ZQhfoUcqE6Ci
DmUpo8ufDZ8ugwLVvFdZmEfHHfAWE6xloXMBjOic5MFebee05ul8o8dZGlSeK99v
40TOKITBaH5lGxr+lBBu399C1kjfehLVW+FKCCQcNxRHpQfvR7kAv96MeCBwiIsO
BQvrQ05UP+Nwk8JWIwMFCkG4XhTW9ilNVOaLw4X8r2aR3H/XVfGsvciBr1IQ1WXY
8IgkntS7jnKMQqHFPk0lAJFvEFCHV5aEvkpI4cXL0NUZS3bjVumG3NfdA8XZ8SJ8
1x3Q9Mc/hZA8TypZWp0C7zEJJbyVSLDA9yptb9yqJPE0KQy1I/49wBsxmEOCIgK1
rveJshtmFRWsZnNZrctsWZgoYShtCnkd03VgZsG5wyUbBT1GjgTm9ugTUfO+xMtZ
lAd/SYqURiPps7SchzLoUNBaiLyF7C2fi6vXvJTcFd17w/sTNTPO5vDX2KyfMsWj
bPWJnz+oG4aDOW3Bcp7FgMqIzF55x5j5eZAUwOtgEfTIiKxHaUO3KGOhgM95X+zv
QrfV1yK5o6HMq64l/8oWrEcS0+ImINkvd4dnCC2XAni9w/yrNkieWbf2/NfSBY1u
rnG6dQ7m8rs1t/pGSKx/ulMi9ry++Suj+Ui+M/mbasrrtiZTm2elIZ9hdUmRnciI
NbZWpFyjM6Q/OnYlxsjeOBYSVX6Ea14iWlUJxrDdSNiaRtAJjvh3FA1aMSZD7MmB
fwt/jnH+7x/wcxeSRsVrmOod2nUv9PyIIaTLUFf1sFgX3DwD0XIhPa50OW+5gTEN
B/jkqxLX0WfAEyMIUtQOYHPrCPvGzi9S+wUmMATDf2t3Sj4Yp3cJckrOUKFqq0RX
75S5Oiqun/DqsnU1tZjMXHsx8QLj1Pt4d4bP+5/d3fPdFpHIb+ZcsCvibmoYv6+8
pxJ+e2H7qspRKDCKVJJmpaidxil+HEM5aV0/vkCN6MT/mpPUEdCwwVAQuXBy3Qq3
GLubdMUmjy8tfsWyXbwUq/pAtkcFUq89tU1zCnlF/9iwkejqOjSvWr+YMEk1xFQS
ljIhZcHrfZLHbTWUbAd1Ga4gCRfEPTDr3E+A2QBgpb9mbH+amWxwLM+/JWNWFUPC
iIQdZWBTPERZJJBPYbesitZSkSWp5Jw7VRgpas4ZNX7bNuBzmyXo0x4dyDpTvMCD
qFDxDTFI+JjgHyaWTdgNtcCORppY1CPuZ+4ndNwsYBevA5LdCJoEdg9GZ1C+2S6b
W0U+4Pqm4XrjhoDX9ICWs9uEGd9iNPKHqUqVraF82oVWFCn9dZYm7tUQhVPJWTBp
gAfnPlVaogVeVy+k/rI2z28OUq9G3ksM8wHbk6JWsABJZJbl/wiW3zoDrjz9+jd/
pz3asRHqpCjZQpGCbo51vlYcu9d0hRaO/WngbJbvC5PI6ZzHy4wWINgLHilKnIfo
TbVSxv0Kbcyql6NDJlWtrnBhhS6w3UWSLrXMzJBOSuTk8RgHZdUQpeJ8DQhOumCe
93eI/9Qy0PCi6ThHX/sjA5R8/aPY8NO5cetRmOha7IjPlM6r9ONZZzOz9pztWuWI
gX0dtXwpA3EmA30x6C4t/PXo3TxjOZi4x5KCT7LYUB0wRIyNdOT6egc8a2sNscVx
R0YJrBnCs12F+EoaSzOPUMlnMs8YpnLd7VkCdgXYzKBPRZgSKruNV+4rxcqRIu5j
yafg8+ITt7hNVoTRt2PlXmldJ36hxGiqcd3xu9fGUV/mEk9w4mQOddqh4nRDvwaq
/p7rSxbS5+5YN+AFhVbsq2Au8ywqn/UFyLI9na91hzhh1nO621wC2JYOhPxiC1JT
aV8w6ejHbrPN7BZ2dU1XkpwKFvP/4/9Ve5T5mOw4aoVH0yNXZLmvJUcQ60/m0kma
vL8YtrtmGuSPNluL1nUvSsY0BIZZGhDXJc+Rg0iGvuUX5lnvN0WZp7Z0JyZmLcY0
+ScLn+AWhKz0t8Oo866wPNd/JeyeDgl2scNOzT/DzE8qo85sW+Jblx18kCizkH49
UlhmTow9Tgg++KZUQqCatA7ATQN2haTabsAp1OCDVd7n2WP2GEh/1tZTO7HwETMz
KtG5C+kkyZCYZk2HJAAmD6ZQR8SVyicdnSXWlYiX+W5Wtg3hitqA1Nj2Jbvib9oT
KOD3KJcUuJVTrZZR/IIDaNCAVs6O/dePZn1tgFYg8UO5Osu4AzyEpa2MxcZ7nMJg
cmYRA+vZFW6Jacy1gCFAYYbDNKFFuF9svWJMcCkamFDXvQYAbXQJkh91RBhVxvpQ
LlYTvFrEnDMmNfrTTgd9HmC+oljLir7UfvgQ7dRh86ZcJl8YONLhu26GVaAzgxE5
ty0hKC0geA2O6KLOt2HXQTiAckL7OXMJcfsfZp661PONLQ9Q1Y8zDWyIUggayt8/
mJxZs8ciC5MEmJiNDxHb76swlOwDNG1N3I4NWwxqrO+lw4eomjWlBtcIrsq1npxn
RmJMM0zDfD9sbeD6o6OGF6qD2Na9pz6IHy6erwzCyU0vgw4FY+0dJa/rLvtg5P/o
qP2xDhYqftdlqHzXn/wKh082pbs7Ok7lRWpU4tgnXi1XhpUiVlKI9SKfOha6HWiM
693g0ajE74uP7UGlrB6ygFkqNsiAb0x9RuzYVds085AGijzqgvAWbxK/orKOMaaR
xhBv0eaH3WulmHrsRiRU/5ANwdG5MWXonEZHaKyFqipbsIoNwLDfGgBCoRbC4071
S4EOYpbtvHZlGjBzpA8sDX3Z7P7UfpjNaHfqV6kPV0HDwKdE31I+0TJE/gHIDm7l
yuM7ez9FNfuYWd5tcBxakY7JcZAfxKbW/901lbDr4G3CEoQC4sYF/ncuvtBJd8uR
w8t9QRhZHYazi8iWThgiugthKzZEJUdEuYbYGpbT8b43HL4+N/ZVz+UO8ywH9jWT
Dc4Oh5K9z9UNe9++Fy561BWu8b78d1TQe9agIz2umPuqU/5H+/f2dPIeI+Dykrq1
+sUct4rJRFTf3mzBkeG0RJPiMIJDhKXVlNKzNIjuc4i/EG8E5oFBbyyBiJqeJs0Q
UrqywdwRrhH/KmDKJsDHkEIPQ4s3hDZJWiS+JEBMHnkExTCf7mpuGvwcl2LgNVZA
ynuxzonT4XZEWOpz83c7a2P+RYDiN7HL1d2A3G0G7v5IzsWFUJp84jSbHmD3cuDp
oL41T2+PhluGgnTxlGdc8eYKI6q7nmx6Xn5w7hPWGlqDh/vDXj1maPmpDhxbFo6R
cqyh/LMat4EHx0lGKFvGa4OaieP36vFI6Snpv700f5/oTK5d+KKiGb/jU8k8TP6U
WUJknz6MB751+hC2ig1l8TPQbUF2RIBdDR0v5Cn5AzFcz1cD7sCVm9/yxuT1EDcx
yUW02PMZ5kmxCf4tHDAjM9fMIKAbQxiR98QpJWBu5xO7NOBQ6FIagbovHAVPdjL2
v1Gp7PK1H2xHh6277zN9IJD75+hA3NEY6QFnxyj5Batvi6185rQHvpksW8hdST6M
QOcriqiNNc5ZrMQuGZeyh7vLUc0nRT00/ZzeYy2SGqjLnYcJgkAVPLSLOcEf7S6u
Aa1t7kZS9Opz4tiGTPflkcXA/2+jqD1xvZv/MJVl1y3lqsMpu/gjYUXXahSZmV36
idkngCRZ8tS/ultS1S+EQABagSTJkbFROOJxe7hRBf2xVwMq2pLHAdSHT5IC+ty/
zZOqn/YQkmY6V6KR2RU0mvWBVZiYb1QKeSCxXGlvJc5D5/sdhn/dfqtgsRBkUz0r
F2E6UHcTLyfHrXFFL13u+2F35PCVGT2JRwhyO2Sc3BW9bZq364C8v4cBE0b8Z50f
NJza3Q+d0zyp/w/YfJtG+lmOBmWlHVQ8eezia/l8w/EK8oBezWfJc4lxgvBnEtIW
CaPt6s1lig9+3qy00mHj7RisacLMPERzTTDrufjJj0+LzTu+PdTlWt9rjingY1NM
YsQktY3tXIePXWXJlRJuV415m2fU2I/T+58bpo6XqWGbj+NxquQOEl4aio8uyXvu
GEcUZrciontIvD5OHo4iQKYxryejM/AdorWlZGoeGt/GCF4aAgDBu+G8j2MnuJ1Z
efKeefLjdALO9aylPkVT1pUPLyZiphtvDbzcq5QhUogCbyyrFd9clROhnJuQhAMb
ZDmUi6dGYjXsN9lt8mrdkDlstcL9RyqLy6n/LK1faUikuJHPfrU77gUneYVGu0eC
ugjGho1Dhke6Rq/K42Fslywm8/wkJOhcUvitzHGW6Us9l1KkhifvebV/wVwbIqf6
KavHWWlza8L3+3LV7//bFfu22qBkcwNIdqDHkuUTW9r7j8g3oiwdcdDZXM7lTeZx
QpsxIDV8l/9oPluk91uKJKlwW+b7SFKpapBv9AHxwmlzMVjZOSRUroB0M4cOfo48
oe6VRy6p0XTDhR65/1az5bR9V3+zzF0OKGj0as8uMbqYCvTJbShbe0Rpg+wyKXvf
aVwxlUmcJo/CZcOf7fzAkHs3uYy3kJxcSprvZ9ouPvMJQ+3bWHIhMPoFCUyTZ8Np
zaAfO2GpsvpIMVjnVpht4JLQFffAvXKfRAftbDK7W9NmXYGXvsog9hpgHYyNDqKw
pxzm/IOEAlByGoTPqwo6xl0DDytBnfn4ixqr0LuxFylKTidG/1mz23LAPdB9e0Uf
cnRL5YuYzJDYDypWletpS2GyihpFxQw3lpd85DMwxAZFiVbbJzk57HB4gHItGTxQ
nPKnqTSTrNQz19Ck7kVq2t+CpbRnqluPtNkbhk5tUroNgBPNvmbyYYXTs4GgFwYa
Oa+wCQ4ApM793ceIMuY0TusJsJkrWl9fod5tvWq92suO71IyC8ASkxjvux2D0/9i
VavlhAFKfdYrRkVdgu9jc3HanmavUgCdgB6lPsqEVjwW/oIriAD9P7Tlo0BX3Ir5
zEgl9KbJ1yVee8lyehtPFtAtBMg2HpDhLqKU5MJsPD3tGc7mamMiLWTrBR3kn+2V
vSaCBQ8ei1cIGzHLPRvvkCG7cRduEmjWpcgv3YKVweMbfL5RLmPNPv9Fk9VgvZqX
qWv5o5g3UJNrS3ZF8zYvU+leGaL+bEoPuxYu77LeRVrITpZbchTm5jvjbsjPRrkX
k80eeLuv+7XlD3ilxoQwcrzUg62YXwm5COOBab8l66mqQxf/z5fMAmKSp9+6dj1d
Ik6oC0G5O0pSCDAkQwNXb6BekoB7xR//Ut3Ht29+16MMPmbSoRE6LcRTKn0Koflm
lIyxVGwP3f/hWF4C8Rr7ftVrIKInCCFqKwTpcZvBwOR/xKrUfGKwvuU9wKK/ICh1
mWrGe+pYwH0YuS2MMNXNwGWZRULMIw0n4zWhtXmE3SyK7v9W5UlRHlMFTaHjtiDv
eaCmV0FsotRqKTP49lncYlXSEF379PrxSbZyLM7WGq39bgLbRXdYVZJ0pim+xHT8
rbi1+ZDEoSHfDJ2oyRue/GsCky/h0TJtdrNtbcxhFMzTiIkgTfx7Blpg17/43fRb
mHkZBoD6lcqZ6zdXjIfv/hf2rpeTe52VsSUegLzR9DLJxTL1RE5WgKB8JtaIYTTX
UEzJbxVuKeB1KZ8u3ePfiKIQ//x2gKIuAZQczWf7nKMf1LYCPgDT6cusfZ+GsPpl
SSCVgl2oblNzL7rrPEXsAto/V0O4IbCtObbNquZBRXG4hpdNYWj4yj1hjAz+Hr7T
Dn6orpGjQ7P05yxA0g4WzqFHiNwPSZeGJQrHUnoD8sbKuFXAAD6fYQ5xRzXQNhXq
itoSMdZ+oF6A5q7gnJ6SijeVETxwV1x51Vv2HFEc6u9I8AxhbfmhVPT0r6ukjA+D
aP/UU5SNffXIx4kbA3MWYrOK2uvR0seLCCUMpkj5TghH/lUp4xxhbJPb13x23L/n
1mnDbSCZAWcKC90FUfBKjMjSGaBe94Zzg1BsgEvDoFnniK1jXBHdXzGr1n3k3jDh
FwqOgdBXkeKFsos3YO+9DSMMTsirwvnhj/IvIrEQPJi6TlyrwUeUUbsCkRgmAgC4
v/mMDjZYQru33sftxN7HnUldoLwthmoOAbqxzB0SRIku5s7NJAG/2mmqc8HU3cu0
kc2gz6iNBEx9W1scdZbyOVu6wmf6uG/VQzPTS4J450RSNPKZ4EDxjvodv04nuq8J
IUW835pwXGP/7/GuEWn0AEsYhDNcIBrP8v+npHymMQpV9nyu3WlpD6tstQ5PkHKi
CbOkgim2MtNZXTL57GEyYgRAWFfdaNgv/zaKtwxp8eauh7qocgWOk9dSfl+KMwiP
tkHpQOdr1sBbeBtvIEfKV4I0mVyGsZsX+RWLKdIeZjplRIfLvfm1A8ov5olqdD5o
9cv3Ydk3/YeijVzak1LGxv6UIpS4sRkAXHkjieOjlk7DJ4P5tMQcF6qXt9Ifw2fs
oCYW2VZaM3IUf28fF3U+fe1lBvygis9MhLUb2VUxo7fBntoJ/OZD/yLhXTvT1ITq
R5vvTVACbk/F2xxRo6mgn45LHGS6rTCKYyNZXj/xCMKueFVvdtUhQTX0pxA0jnOR
dpgtrTcpOFM5hi6WwtdH0VVcTdKadG4C+aMMDoDVIPPAtCTfejdkb2IpImtQas8U
VzB9J99juUGz1VxWysGmPvHtNWob1SR/2n/S1abW4TEH9K+NTVt0DuYxvkoeyUps
tPnGgzb7nK/Wu6qscZWpVIoq6jESjPRJU9lm1Mmw4qTpruqbWigL/w2QfzJ2xBWT
A/tt9SbvbVxJ08zqymjwT4G4k8qxngfBFlvD1h7aU3Qqxhu16VRFrUoQNaZI80py
9Q5+syPFztMeOhAaFXCNj2AXKnvwZUnAMs5tepnrVhahjo4aVfVIWkaNwaqHzU6s
9EFc3eN84Uyxjo3xCQrBaRlgN7ke6lTyvHXjuF46u/mmp8lsy7RDS9fuu4dpAYvz
TWqU3V0eSX445L3MnCu8TxZQABL3XG5ilPvvFP6+PQon2gN6EC/O2JJCW8BJTQL7
yi339N+wnyhLQ/H3fCTST4PbY42O072Ot3ON7e46sSw4lYsALqvO+sYZMKqZ6ZsZ
jBiiyHRH/qrm+tqkM9aKnK7YoqmNOP9fn8R1jEWN0koRJhsrXPUw4hiMh1Myb4oq
KpLmjUtcBkgJiqrPBo6lUMwiDyjW4kox/ff+X9gx+gcTwIbpnPVpfN/hHC/XQ4Gr
/paf2dqwAoPScrwXU4TdzXsbnXPl7Nab6bYzHRcI0o1SvUsuFcluAUkYuk3c1o21
mtScg7R+iWVEEqRzZzvvovfybEqcxCgaqxHJOLod3K0z0BelNd0Oj95Imm62PY1c
o+scilK0xISZGw0uVK93ZTh6Q1+G5OABV/uusRbt1Hgi4WgvIs+PIHFnmdONtlpW
KCOU+fOgWI8vyqdWV9/polLuSGeaWtgNvP2bVSD00wR1gq8ZrB/pIw8apcbLqwcL
mKqy9/XLEzVH/g7ozQmA6tztNHAB57BAJ20jPhtBAUv6WWmQ6uN+wD/+d7A6MCnF
BkNll2CHyC5IiPSqw1gH59yZz34WNzH+P2tjF3vqWQKO5hGJQoqrsJUtBWhn1C6e
iSaYHZeyavJvSoW+INkduV8lvLq5UVnk0cyRol5GyeMFDr7qOGO8/Oes7IUSsZT2
FjWo2zg7cR18WdEx8HyU8dbKd5j9d2Mq9E+XmVOaLCUuiLWYvuWcATLyvA9TnCAi
zJ7a07A+ycmhjnnAdiIZSihnUPzBIw5FzJH1pLfP6VyDYuqZe6M8moTSIullxEFp
/2To5HXUsRpUPg2yvhHJYpovlmmuV6J6U/TRLqvgfxBpIhO19jYvWhQb1sLB2N5Z
wfUPOmZW1iF/ngxSm6j+q5wz0uBNjQF3icasvV57b+SfRamZykSjtnlrGN7uHWqo
rQICFfY6zEDcW1U+2W2erdrxx7KhfrZg3cD/F6U/p8DkabhhMet85Bmns0j6TqYO
0I3B9GdMK5DVMpv7IVuz7krD1OP4srZF/vVk55xCVRUcMlOwUePwer28oc5/gRfi
hVozm7sj4bgjFrPwQkXpTPDrCjk//NKzIpCwiGkAZA+xG9kZePrmCWl+IeENV1fK
+SbnI8yQQGujSk0tLTSKuq+hZOtHLmgZ5QBeD12dvC88NBOpbNXZzNQDB/Wjjgi9
+xIo1f80Ao8A/SDaWt1T60GdKVfHS0S73eYFuMcGNdrUBEHEvLA0mWDFd8ulO3vh
HAFPQIZcNHw/fdT5TamvMOVfN30LGwo1Ff9uzSzsUtzdoBFKW/pQKlZKUYOEBf6w
76PKNlCObpByAzkg0BfCqdb/XZZrOAmB0R02w0Fa2goRh79ITTc+c/l9Pplerx4/
WKhZDbyxEP8+UWzmlT2+GK+bqcerCsgI5US1loBKdWzE4hLgVhmPh6GdbCtaiqFZ
7KbDlMBJp81xHKPfG9wQ8NtO/CQ+BA3ztrvCdlFfneGAAgUqdDjlorTaPVipBrTe
qu72mMzCMOvoW3eToLdLUEPpobF9mb9AG/TXpMLBe3DeAGxagO5Ti0jPWR7vK0R+
dS6Zp06CHHfSh1NyyeTiawWrNmwV1e1kxMQll8hoJ/D0HGxrLKRaEaiNzE5n+4kZ
iyMqFesQ9qsR4T7FycXQQaisdcKg8nNBpgmToaJsqcTdOnhBf+84+bPu0ZNBkoPw
Gs9zREbG17t0psw7Dkr+mBEowmY14PC2MWbaBnMDOREMXHVQfstRnBMhxa0DkVzs
DOLL1SB1KLHf8hxfToQ8oD34CLiAsj/XL1lIn3O8GcJOE5/AOtKJC1orTTxr75Xj
uFZ+UJDBx2Rq7VwcTW9tiV5C0XW9Z3Khn/QtSD6DTJr3KJkol/gIcitLAX651cB9
lGHH/+/vV+L4wu+kaM1pUdm15ooZkGGLXKynCE1yMUQlqzRp5CCsRQ2k9BPlJDcH
IzwZzlitY9PGmQBmF26OZyCkCI7fyEfO9mm6MYnYeBXzXL5fn2NoomjSe6TB8LIg
E2anSVxu9wT3Dvhhcmb8WPz3ZOzki77H3wYE/N5EOqoHC5y/MRBhGo5IzydJtvJ+
SLnHIz+eF87D/R6Z617Y0iuS/PPXEsDL1jieHrjK0IfmAtN5N/EVI4zaaD8K0TYe
u6zuF8CCX3214Pc/nKl8uNTQaw/jVxR7tsIStgqrXYfVuc4cYnYFsHPfXc94bO70
Mt9YmMMdfNfi1BXkLwL4O+LX5Ie/xqcluOOhxNHf+mx4NGb9aMBmDyPJmN20f9p8
PBYttqacaf0UFSPgC/qLilB8mU19BDi+eyWaeGtAyjkb4aYCuKA5C41dLYBX9Iwd
aVR/d2BNpfc/xQJws1XBjrWaau4CVxcNh+hF4GqQivCVolWF9kiDrb4+VobNuZtx
/PQw97LLz24/p2qN6kGFnXo+gTZKsADu+NcBVpEEace3fJeBWu3GVDJyLiTq/tOt
9wmcE+gkeuw0tFvu2i9zTqnO5XzwtncJ+ohqygMQkfLeH+WTZu+EGxOQ9xGbbOfy
poaZRltZh4i8EFXzoFDV7eHVAm3Wd08zd37SHlPVNjou0TDG13SSRmL+Siv6TywI
D91Qq/gNTCfKHPjPPx1XC9aXuQVVWhg1zjZzCk3l0WTPljvWuYKXOB9h90iHtlAI
e+yXedMfb239K/IEqrrJimnd8G14d41sOzjkvei3Zbbmfc81VzVHOtPWot+0x26R
3659wgG0T4Cp6EsBZXdZUHbTVxHiJJzlm/KuJCb1BybFqgdyacF0BnfNSHY5qd/A
pZMsAr+0/XQ+rOWyk0KPx6/Sa2LmizmxcuvZoIRvQJSyN3xJs7c4lCIkJ33XGaJF
xBFQgOzmIyRJJA5sfQlgPG2akX7weCcm0uFhior6NJNS6cp7E3w7fo8Amz+xoBST
4QSXMPe0prZPaZ3aHQPonBt95Ub8gNuUFVSy5Y33tr+IFeTXJqoeWikyNN1uENN5
DfyAZIUFUyA17q7F0d/ckh8pLGdclOPvj3uxu2mWsGmWA/kOTTAmXN3KpPEZi7Ay
Z2rY/d4qFYqMgW7TXrnv7aI78N+Gi3aaaNnsCVjcixTj+nX5BE+EFCj579CgTxYq
k6/cQIPiL2DwkA3QtnsGzSLhxFjsnfNf2PoMvpC8vH7ObQXqJZ84mRW9WTUeYgAd
mwUfZfdt1oL6Oeq/EVLSaGCyhCqPV6skkjf3Q2j74PM55vptYZ8dU3u6B7Qfpq+i
Nl4KexbJWJDsvZmMZMMvYEW9Lb48+ORAMPNaAJT14htLXw7qx0N4eoohOgUwIndP
ME0/OX6ea3pjNcRAfA+2bZEw85UAjyVCqT8iMWyIRPzgAfcS4VI1Gubhj1ivhFb6
l/MhNSbGx+qZtWXLIu2Eu6q3dmPi7GRvNlNutXlGzTJ6J7vV+fUziAptScJ34XOo
WSJLLvhXnuK8LvS/B7IGMCwKbDlVG1xbgPNKlAXBa1YWt3+kpHRp3NGOYklcYtaW
0JpPMkbet3xjBf1dRN9jE+OAoKmbaMOq4IppXN/3XiqKHKRG/yPb7nMUZLM486qR
BWzDty5oFbDdPgOiZxBIKLwAYv7BxJ8Yf6x1LX5IrfcJgM5Fei3SuyLnpIY+g2b5
53qipBfuM13eAg6CkOutqaWXsRngjPXuSoyb3K0N8HxHFJWSrTBCVqT4X4bbFFWa
Y0NL2IvIIbekq9YMfnx56xD95MmKS2dOXqDi5agCCJO8V3FmjkavgUyYJNDO6VSa
QBsMPjL9e9RBFOxEbpJ2uPH47aj0q7FHzKaZsHDt6W0TY5ErxwrnvcRfCiNy13N6
1nVfTIOlHYDOqvjPskdUovtXtX19KhRinrFWYmd6tehPdF5f/T2eRc9x6POpuaJy
bulqOV31ktqnjmu/hecNGkJ9ldSMySJvundZwL76FkmAZpd6x6PHP/D/cODnuh/p
hs9UKlysa6S3iaXsb5qxiOve4ZacjWYtoZXBvHSaNwk87mdqxBzk0rmaJq6QXwcn
Bl82k513YIzHAyRSg6SrHhhKSdzCJCZXfcotGqH1YmKq/GH8C5eePgBEtQ41gzjW
cyNgfZ8W7lDOyLOgl+z4JHdcFjFvMTvmRi9uTB2R9cTEc4neESaVfV1/kny2NoIv
QVLor/+ThHzB+dcm2fyAAHSPy4OaMAaQMtmjUxsz/vnNAQE8+9ccU5UwKrgaRAWD
2ML6MFOo//IiaaVtZdZEIqjESmabhU2bHV/xgq4+GeoW7OTSQ787Wq5VJO5iuNnd
S2lS9F0moXWESG/umtI8ahHc0VwSugNX78ns45c8MsC9614vj/nGw9uHYlTAVngf
OBz6F6t/xU2LzNpzRCM0DvOHi8NIblVgRkrW9AYfy75VsblanacnwV9bKwkbBClC
JZYmteX/URCchrcAL5Bv7wHhYxfu69bLGAqCvnq1zcRx2blG4RMuSw//0N8otjaz
r1zWNXCZMCBS9EdB4+NDtsX41+RHIjs8mt6Q1yjTlwZGRHpfn5t48LW+ezgskyk5
S+zdhDyHaC8sfOcIuV6Y0iWWKYbwIR2ZcwHfhJrEoS0R/2rB0u8O3eE55qLKRC1k
UAu98AXJkB71OIOj3bniyr8natKDlEP4xqCLqz484UJWciNYo3NdhyvXRSCx9kjF
jM5dQXx9g3E20Z+FF4BzMtGhDtwG5JTuWonK8Qm3J9N42mcpwb7sNYvBrNDipROK
Xt8W+9w1v/paf9sO8QpvJw8uuV0Q8sn0+C3ESBEgCQVVn9YHsZiFiL1qFlqlqYH4
CKyFF1c3JFoGWdsijckfjaGV7IaLsCiOKyKr0gJkTpIkhHc13/K5rlG/Xx6K7R/I
674dFHxrrhInT6EDKpOCD7SrJkFArT3fRmJlysvh/GJOTb2Vs3tZkY34djsA/ezd
f92b5Yc4JaFnzIJtXazU45Jo+eSObq8m7XT0isIE4xr7Mh1sJ/TZy9/QYi6svs09
FEX+vk6H/Oin3EWrB/SJeK7phKS/KqWAtBEWu0BQLFCR4fkKNbZXg5WnAjEnX4CW
3tV3ExltadTeJl0n9s24AVLHvP7PQgfmCjT8B/oe3+BBPEPf1dGRBRe/CfBJ1K5h
bFMCl4bXbpK3C6cBCDa3AgRG9SVVhJRK1qIsID1lT9phHgW05DSssKK2+j8CWAOp
sWUtkGH52kbKKWdvfUot0P1zxK9Fxr6eiTeTq+Pvn01cSUYWp77PG8QIEaa+ku5Y
WKyfW8ahcXdOCWT0mCvvtf10WQ63ni8VF/C1KLo9+5VTX1jjUTXU4Hnih1D88g6b
3qBXTKjPWTgRjSodtGtRHaz9yztAeyCEPRKjgDX46oZk8hWw2bN7KRgrrb8ljKMk
U4R9BBUZM8KHzDR/pWB/S2yPhCe9VgexG2cMxRhnfos/LyNWRuZhKivUkLpsm+oZ
0oiGRG9cSxLvhzkQf0oODdzZYOHgEEX27kRMnVCJiePMP0/19NuJ13RCLTR7HCqW
Z+rYJ8uYX6Ob+aAfjazlakwpHE57r6NWGLBFNXF78ZRHP0EvUR9nTLzYpJZs6mop
No93JJPjFrSE+C6KHDSACpctCW7RkqaF/X/rnL/XhXWUILCdDAcxfkWG9rwpoaZo
rmoLvJZ+k7CZD4TDQZqtUqa24HhWFKgbcGmXQHd7b05JBHgQnT3syUJST7Lvt57+
kKCTQF/8I+TiEPdQ01wemnri4CvqAPTx66FwXP2edmFiX8b+90FU9x/2Jpve4qxj
CvFkKDAlGJcc7CZSet7PyWLPWhbDl4qrvnf9oob9KQuYWqJ/3BayiyXVKyT1G9fV
AjHrUc93LnXOzP2p+iU8t07LWidb9OcsqnYl54A6pooiwbGtzGlq1D3yQQnbzCKY
ds2rqCvCF57uwFnf4uwHSJ6lirE12hMN7S5EgypNPhbKLtlLU8KYSro0eGbYPKmQ
dZa9COaKHKDoQfXLXIYsXay35Z6SHHk9kUjhr1rljKB5c339y64miK95iN+MEA1L
z09oOlRavJYnBbR+dyCGpMIgXh2Z3fOI83kGcQWyE494piwNW9IM12hosbQ9RqkW
dE1V3Xf8e6hTPQTuzz5pBf412W4+8C0phhUv+mf3mrFvIFETiaHG+z2aZ1M/c2Ic
fjXopvl8fgwa7IQWAOstmYmitcZAvl08Vv1fxio8c3D3P4AiagF6KA3vvjiUe9+L
aIYvcK0kEkRY58XgMFlyEXfyUanbnsHH4BI8QjfgchpL78wSDghwzGdQlOhh5yBQ
v+FtJXZatzUjgR3PO5PzyZ9pjY9HVTSVx4HjNHcNpjn7Qyniz78mWLPqhSc45lbv
rbfmvXQm4JgYu5fNNl0D2t36jIJ7JBEz+XH6CTpD6sOFpOYy8W1oMulNAo7AXg4E
i0vJndZNfd0PbAoegyHJPxd7gHELJ1XrjGOYDQrz+WJ3vupi3YdTlapLbLLeQJUu
lQQgvdXOKvv2ksWzqWvzBIXdJKPzzBYnj36eiJ006bM+OhDs5l9tb1h5gebSC3GB
gUFCT8sAAlPOiffHupKHUPz2hESp7T4Vt1PhFuPUYA+kG4hXI41eLhe4qzq1yxgP
QqmgCu5LZztcwO1DJLNoZWHtsSkGUj1oOwgEO7cWDWkY8d7uOr5dGB+aB/nS3Oi5
QQxwxdhuEUMaRg3pYJjWZ8+9MY7K+1YuKo+0BoRu0pBowZyaYeRRKsHa932N4IV5
1JHZvfvTXFZd4B3XE+xMg9KbvNZzIQmQ3RajPQ2h0qiwbI7YupL6saDHFu2S9HyR
WUzVmPj5TxBd2nTatTviF+CiRmn5k28fRBPc62we14h3dMq0F9F/iKESHpUbDaEg
FzdRW5ZJnXPi07mN8sRxtYYy+LPkBsNmfNXx6zAD/0t/pArNj99WqAYkXlypjAqI
NTSI+6bizgUNMMLeTLbInijUE4eHJzXzSbiItmGleGS78xpVacBTxiJ0nVLVyFkG
0g56RvOuY9pIfqHBeqCQPoiUIaIsUwSTNmHqdozWYGuvzlZshwfT0VrxuVkSymbQ
pP5h1HHDFE5zL9FUGbHzCP/mga5N3Mvki9vTvnStApeKVZ+5v8DF5lntw6BAFRK7
bq9jZc1V3A7XT9Zm/oYJPj69ZS/MypCNxZeRdBBWW1FrEUzwfFXHOn9iososFHtt
bYKNxmXnPS8Aki2oP0KJ0isH2Py2+/4rkbMjLB1tWNq8lEFXhyHfYC8UobYDQ4vh
qBiGcPkSq9fr/Ne9ZnudIOiCLFwQvuMKXWY154S29Rg9QBSC7FieiwRUVS/4dHNp
EMjzpWR9CyTrKRMCEw5frLnDeANI/QG9EYg6QEBI9p2uG1wXsPOH3tj/Fm0HFPgo
IynA/VwYil+a5g+lwEw2l1mYPIyenInlnaivNHh50gLNWz/+pLBF+YKvP1vb4qxE
DHxPmk8YfOcASAlN/TJyvSXKbxi2ZBOrrqX9fNyolIB8rzcmsP+Cf0gwlBCbW9Cu
zKE9n/7Eax0dANEUKvHL4HDbIsiW3+CVxZWy7JHT+z05WQkhyVlTDGpY3tt7O7WX
BMhP764Qcf4ZcThUZVqRfChiFTXwmwJZ59jUyZY0SdFovzpMaEvpdb1MQCYlMwCC
17yvJsEK+pRY8xPe+bzf+mD3TLaQwa+CMJgGSPdymU4gjOtaJDdojyi+RGu6JGyC
EI0EL5zLcn3I14F9XLIweNDkc0UjF+X8ubx0hminsb8DO57MlCt7TNaN1FxkGzSF
uz8CUlAvZYMomdWgoAmbwJBLUGaXiwy3e/BeXauAUGleHf8hx2cUhdemmvehS22v
E66GQkokDxbGv1H/U5YwlF0oJ8QeBOM1WuXdy18jSA7RYqde/eBmTK4WlM2wZK7W
JT/3DGAV9rYFUBJ06qyZKUvWTDXU8D1mOGGZCXTMSG184zkv4S00D0b8i0e3B2pd
YIT5mGvKjbNvMwj3gKFrJLYkyoY9DM+vwcvdz07qZbiOSuYkKzWYuVhPq0vqK+o3
Myu2ofQcOh7bk/Bygy4Sgt/d1U3pOHUzCXJcMUu2eHAy4Rl7JN58TDMBjsUIwR5o
PAYQxmhaf/myEtK8Jm2QuHaypgAZYUX9KKUVJs81kF6t7mSCSe9mkQTmp3P0OdbL
lFtsf/bcXPXgwTtPCOxb7M/LMU738bdVEy8b3x79ZWKZerWbrPzct7iCXgdzFgRT
rBS/2Lbs/c3sY0t9qAS2RbhtZ/zZYkLEnCrBDzFWWfQ8KS7on/4lqQWpluWxSr23
o+DorV9fftZJglGXbXlD+etKnhiPNdnEqsTpAiXHrs2eQO02dhIsVEqoeGJsnTvd
rBP9o7WTOKrmJqRzLNBSfaNrna1EnDKit439Q0pX9MFlrJoNr666U/ZaS6ZjPs5o
fp75yUnKJ8yG3W+74AMN6yA9BoD0TICMhxqq3LKsOxO5A9mgoNmVGfdiusfNaTTf
B0KTOSn4rocKiCbvdJ8AKcCj83NzoGQggiLdMxpPh36vCojnf4uqZWSyom9v3aUc
3WZ/RAiZWwBms1CSJp1dFBfabp8bzFeLuFM2blFHnsFfmp2koOBvqPOh/d43Xvjp
ryH6PgqG4PMmVWsuZlVOeETD1pdP+1WIAIgUG4irD9zS8csYjVzs+Xsfa+r9lBJs
CJgKYliSERrPhbFAquuas52xf9H0Vu+h39OfcKFdhzXnkkC/C4TM/bgCIjNN9Kbg
hWlCkX21xqCS2ydYT7316V/tg3JojoVrVRQsuzJSgp2/+BbbW9YSHN3tmXptmrac
lPsbTOex5Bejx49wEjyqGQrQ8yFDkoPQed39pDa+gwY1op4qB2koDWVQuh31lJkC
BtLM49DQbP/VMz1/kcMm1Yvt+jVSPEmiR8LDUYFZl0lI+/gagSby9R3rga46Qar9
Gnac2jeH6toOPlfxF1UpbvT813uozcQboScspEQEdpKnXVqa6npR+2hTmG3JkSrc
qFUuqdjQFYc52WpbvHwXg76WcTyox6z4xvp5hzNC6ZiodHPeTQ1GRbMM1ECCvH2h
NJAWxYAkjaFV7p8iUtM0SSOJGvo1m6xeqKd3Wfhqez2B0K+S0+Df1PiJkZIMKCRN
iVqjumpMrX1A8GaI9bRHGyXi6iuAELyNish7pJxAEviJnI97737d+SuIXyt+7sbr
r8QGU4mMr9yhN+UnhXekQ2LpZ7QIUX3IQC7Hnt1v864RiFi/5lecvFVj8A1G93sd
MEjRpIN7SLQOkM1rTcBF/2tpXh7uXkYqP16x9BDNxQeGxxyrHbCvd9jWdii+MAbC
7k9BVvvkGCYfzd5COiVdTf+TAZPpHvXAbg1ris5FA5Rq9QNTXVNpcg0YygKxK8tx
9ge8rxNzIBYp10fziP3oq+Cj6Snfq7uzdKF8jQ3eIpMl4mtaxLC9yVsmplOvb4g/
iHfjUknzV3sjMQACYII+tNJPI5Vds53A5NulmKiU6I4FZ2GKbF0ykowf3E4JqoxQ
HrAd/SafI7tN7ZHy2ECnc1G2DnRygDcjHCYr8e4YnkFBr1tfhujVlX1AyVUPCP8y
00FzTRvaWUI39Fu64EKiy04suw/PtQiFdR23DMll8lNKOtkOlnSlfRjLyDxmgbH6
PJ/MJzhbizjXloa1Ut827Ox2LqXYKSAJongtIrygc0bAPcNo2jOC5ifm4m5TzPeq
k/ixJ3MJLwJku4Hf/Z69W56mQA/KCCndg4PJxhVl5Cxt5iAMNMRHhsnNQ7p6IRxS
mwRJufHWah1adaU7ZtTud8qb2+meLwLnWfSSC71z4YMyR22fJxG+wlfyM+gVL71/
MCHVYcJixlXdEzN9iMIQUtojcqM7GlvBDX+Qwe/qWDxEJsokkfaZPy2rMYYqbtR6
KXj5pW5E4/qEXs7uSI19yaFBcUyJ6ham10bRZsGxFVvYmx8t/KjXQyjhojc8UarJ
jtEGsMBrZQkyyoevd73G/6VPMsCeg5afgq8BQQeSUGICMMWYI0hwxHbn+qW7o7XF
TQrjTr1aBXkK+fZpuD2YmA+TGGdBNmSHtFlOGOkzzwZLtCbZf3xlFp2QgTQupr2+
pbTt7SqIHqdSbD+oEwx9IzK2jkWJip8vzgwlNxxZDNt8xwAg7wa3T53/nVaSqOyw
7SGgw7lL49OBwEQVeSYeLiVjuNAnMZYKJJwlyW9gCWcNZ9Aon2cqMuvA2W2g5oih
OkaD6T5wKzn8xSJNzZIPM1H9Lkzyx+uMAGevIVTVuztdQWzlSOuqzgh+UnaBHGWs
bn1CkCrCuoQMdnk4LfM0aAegiTgPXQGkbX7Crl75wz+gEE2uLAKqLW/tF5DPeEEz
Ne2VauGYJav04bAZPNhVQLR0hABuxlH6evemhWBsXxbrUckvvC8VqyK6+LkooOKM
z+PwPuW9rwV4tRb8RCs7yD22vagc2eiyjLr9thhteAeHKZMdloyNbMwlatkRo0VK
BAu7JyMyotrEP4HCFO3GlId2I3Weygnu+GiS415indacWH1wBqZpfyqTbfEong2s
Krl13G8hFj2Jve0JQr9qkDMPURX67O1xElMceFmnFQtINFFbpdJRxGLq07SPOHoy
t3E4qG2h5abZMMgx2R/l498df/r47SA8UupyanzCo65Hd6Myzh3j84itzjbwMd8A
MBYDIPhOroOY2fjOsQlSfe/ZSDs252eGhJY1kTYYLCpbmRDRUO2e8OHuim3JPJ+r
sDuHQH7ZTKafi9t8NNo4nThESLbYnxBlTdLhfXIdiYHMQ9R298hyCa2nZGx1tvfE
mLkfY6RNy1WCkft4XbAa6Y2UPBC01nm4caYxXXae0uIgk0emGBU+90bx/MgnTcO3
d+OlJUhv/QbWdfYOkQxg5PzS3Dy7RqDTQN2fvzIxC+goOR9MHv4HjaKFOiVaEm43
dag1J/HUEhi43GBybtCUQEyeU5nV9BU1ND3F44vGGdqcE4p3kltBbZEpGipKsarc
bTM2wEh0KvmIyJxddtXQsdnfU7a6vcTC7VP/CyntgNpwZ+UMluKZq1D5uIKaHsdP
d83IMt193vYNPK6d72MWjXmdUIIrxGCCmCXeEU4IaSGWE5Ed6KS15PZK9RJRvoyS
lJManbcaXOy9mIASpwXLQ3lOUcJWQfDoaa7dJoTDy3VH/JY+DOBBUX7wteRY6qjb
+3u2/K/wuRV8BBiFA4dtDRxbj0Tn9lq1pgHu6MctXyW20V6ubf+CuTwUlLNImdFS
pWbVIA2yRm7An32bXYHGQpd9ZnYs1eiFUBRcJS/6gxk2UsWcaGI/qi81yhOBgvWC
5yOe9dpg+F/vYY7u2Ey3gxahqLMCnyFfJrsQ3TrlyqBxh1uvVlwcvUIuL1adF24U
t4aGZqAnFBxQ5j/QcZl/+QaHvAuYu7n7pQNwrOtHbkGk7RS+45Eh/V9Nk0VkFnP5
IVRkBs+ogW4kEriN0O0FDNzSMk3dlFmbIEXLQowjETvWExnUtRz36rYnj9fytPJb
f7bv8SC3HZFRK18uR+IbjAwBYNn47ZJewIgaLRRDvbTA+5rlkSJB6Y7jxkyJuSgQ
ttaw5uy7kUs7cJ7POVUwB+qn3sCeHsobC4dpBkLdfboUaoyJVWyzEFwfWmGIa3NV
LTMUR5VuLo9LWAB2FmCEp+5gx0qy3O4eqQgv+06GXjYgPi1dk7Xn++OvrpzljjFf
mXGeyrTUw3CKNliB2oEKUssO8PK5tNeQ5qCQQAzs6Wqa5mIjR8B6uVo7wLcir4Hx
lMKiqim8TSHc3HIRWX3iKtoO5sDXEBVlXg7mmRsjfNtRDzMHLmzsKcwha/xrVGtS
qNT1E2bXsIP6LjHCH/qLU+IogpIAjMNBwXGiPZerKJUbaHOaZhyN0X6Wmr27T2Qn
c6Y0Z6wCZjbLYBxbYsWg1yPVgv3TJv+eaRLRen7xw4u9O7sRWqBUCK9GqZcK1c1O
sbZLKq4VGIMFtm05fbljYKzVIwcgXTon34vwgIQvfBXNh7pgZHP8KmiBLGagH5M6
25pmSnsHbqQHFK+9n8owStINLvv4kQSr7amLXK57TTnBjGUakYmhBVYyUKNJIwAv
coRVHp+1Qt/EohtVsXfDH/NhoWq2ZBpG8p8+NhFzMS4KTJd36FloY3jGPuXV17+U
4lTRMskjdZKpLXzF7BKDqV6QHiWv4U1QBjL2/Y3VoT315xrhNlKVmkKzALB7TFG2
wvJAb3Fz4GS6+i6f0GTxZQb+exh/p7CzyVt8oDuCWhyofOOD65c3L3Z2CE/p5LfP
iNRfZ6HY+pcgchik51YBFlLddw/1WRxL/sNbOJ4MpzZpjqCtu2d3ZDtyGix0Jw1G
1+JDsdlWXMxud5egm8NBt66mQe2vxx6cCC8gBQsSB2hpig0CfTC85xdkSmG3N2Um
CKy9DK+vZ4GNKW3axyMOHe2LihdIwcKaDhqK2bdwmpdrdVf6PhvBtp0xIClh4Hte
VSsBD6yz+hbeK6uhxz4b+gSuPeRNxv+fzMGJi45+47YOCV2qM6TCfBxEvgxx5NeX
bwcHUmkfuXZ5jq/UhhZzTc2olRLG+Ukh4uu7AVy+rMFnm9XnakSmMQbkXCds6LZD
HeI9Dil1n1u0ufSlMLZuDtuAfFwUELiNlpFkRmVk+wiobMM3PFWdfOG5kxvj9z20
RnMcsAhsDCzxqmSt3ZKqM8qQ31HsSTfBt2ai8pb3NP6VFg4YmXIrQFrMJpUmZ+ty
fgP3ACe+l1q5LZUU1NtgRDTmetcuKOUdMwPF8IeFC5jpPM5DIWUAsLwdag3f5KUb
AchDJCCYz6AohRbiwhvw0IDxs8IWqtK83zLPADiLThEFDp5PoUwrWnZSXVYVQDgO
Cw5jyKcY3UZyt0QetenP/EEl70kP6OFp3+bvFyU8ZdTBWuudQv2W8f5NyOlXMWCD
S7tFeTDp7nLYSL9MeVqum4PTlRnIwnARg1aV9sPWSmoYp3/uzFD85EhfcsMgkYMK
Lr8xDgq1YpQeCooQK1RLGZ/D9GbKQdsuO3dJT11PdiVvGMQFYwNtc59A4JkJ016w
EXZUBOpD9kdp4DcTwtr1S/7Q0x7LYZmWYd7i/Sl5AxHwzTYh/HfNbqQGVGg5bZay
+H1l8gQGj0+lyvKvDCp4SqjMyoDV59rCqwxUmv+b4K+RU3zeJTfGTM5vUncx7fiL
d12p9/ohU2HNDnNkUSZGMj1l+WPohTqfKyadRvIier0+6rMQfaTtcQQuY7RN+ciX
5mUfteZhIqh479vY6PqNy5BYSgDlAWkazNzKGQS4zPvYubHGMXfQtYoQ5P8HGgOK
1+Jpeu3Tn8rd7UK0NcnVANX29N5NscSlfslbflAqpKISDfSOGS39R6g6GMss4AvS
p+gEhNKmSO05r+tGuPsbBkBamfSt9rsKADO8wM/pltuqgiCHX0exMPYO4V/Tjf04
uojm2xla9tVqx39IdUa+zoDxrF7qGLGdZAfMEq+stbp3I/EXUqskZgG7ouqJigTl
lkToD6f9I7/ydGUAghdkRB1TcIGsIqYWHK9gA/Yq/njuMra6Xq7YP+1rdugWMniH
2tWO/Bi0OnsvXiG9gimApR5UGBCEyBGJ0schFhOW5pkLpJkrdCfNVqbIiwbSQlnP
qR/jT7NZg4+y9Ba7FZ5CEoEBLhns7NgvF794w0JQHjTYQpxIinUAFhpXeoF7HgYE
8hVQq1rDtqRFbQEgoyBL97XsuhA5ThmfEQGX3q/JLKax6VdMkAGdRwdZURaighTN
jqJbsgOlKDtl3WH8WQvaRIabh8NAkhZkiN9AhhPtbwB+NyCNl63M/0OQ4VAO644c
Vg+gL8i3aXsRwDdguxRtO2zDOXkmIoEdk32nMkikxiU4SmclZuo2mlZNLNELuRvG
IKBp11jJpyXlI9abqw1AK4p37b13FBwxjm+4jhuk2Zu9ZXgtfceSd4Q5hV8nQ6c/
EGiYlt6azbzFB3L/47hH8328SYF42zrHDYqvtSj3tGvGL+SFosApuTiiu48kO3pQ
OX9vyXXuby6NXUUDZbbOZhq7/2csj4/GNwtOx6sWmnUANkDgmBlAhAaqpEyPh/G/
ICS0E4nCina6ooUXkhjN+pMpJHrdNdWPjlpy2IBTkqdyPHByRLFb+A01u2cKR8mz
fTRasq7+OtE7FmnPvw3UL1XKaPcVQYC7HqFJkmJxTCjUu/oP5fJwFE3fKkQNWlId
0iH7P0aI/4pQW5XKT0bTfvlQMU9HgbBFXaTQJequ2V3Xg+KNNf4R3Ao+IhT7n5E9
X0l5CpbAoNkIuUAi8i/+v6tq/TTYXsbJDA2vStfZPlshowEpt4AjyKdNObcunKHF
FbMzzlNjVyTTG07ejXdOL4oFyTpy46HPOcn7ZNBEQwOA57u37YEafJwrGsKfg6vG
KSacSHO9YjD+/Zjnbbbg+lFNvIgQnck+HI/WA4MhUhyQ6P6Sv9aIpCl4VMDl9Ksj
QVVN91cjRwznTuQI8a38Nuy1sYibm3BxkWn9NgehtafjCRaHy9JCdeG5nQLb1nym
g07aovo4prjvljCKaaplxbxOwcexuj+D9R42EqZCBjCoQt6IipdqdZ656449tosq
HvAVhatq5Uh+ThwZd/dOC5St7qmf3HzrVO9kOF4VzLl/Ei6ytlHKZjZmNgJfN5mb
icOk1bBKPDMrrDlqOfKyJTB6bm8i/AxeqO4whycPaDDoz6qNdA5Y5GLiRZpzjF73
HbPZxlmxvlpfPv6XKyTKfIKCz6aLjLs+0o7YVy5wH2ATNqqlzd6j1h7CdS4k7uO8
TWLhaVIvnv2htoUKGn/vZhM7MgDVB/Ia6ZAzUuVKF8MOGgoIQPj+wm0HegU3lIWE
ABc2ZhDsq6CZ1zvFt4S7V/abrcjDhleNPlQoTdygD90Wr/+9A2fcGbsQ1bj+sMv8
Nq7Q3boOK5exF7OoBfnorUudXRCrfNrfBzNASSbwwlTrwQ0DnKchn7Pg+e/ETS66
Vgj8VCO7auKK0nasl2hhiwp6PVznf7IW2GkiZ61Khov8brHuxWTgaWBwrT+mi5p0
RGCrQGDjVkBEfg0eKCvFg4nezy5egcpQJCBs/xRrN322CmJO8KhKbVT2ism5aAgR
d8sr0bCdN0M0eCwxvgzjFpJOfUOv1PnYu7gQW/AK9TeztzHV5cOJs0qJ8A0k0lrA
Eqs7TEQAKkUA420y31D8KNuxvdub5kjxJK09OOjUNoVEJdW4T6iYJ/0mI+yE9jVx
EiNgUg8fRe2pQRBhJx3+h25F5nt0cZ8SJtmjrO9H8vtdBjZUhSQ3Vj74knUrai7N
Nv+mIFIBqczan5NcmyZ8gr2Y1O6nzbU4ZFmti7yxOt2476d+jrshbEY4uDNLdrbA
QsPt4HxngIc/y8reV2TKHZMfyJOnjPsInfikddPNsCuTw2VGnaBjHWn5ocCy49hm
YFdZeCRoAelpWDd/vT6qSQv8Ez1G+ty/6CiVMrPrYjgFuTqYCvEts6CxJTmz+clw
dHADsMTptdLHF3vrr7oMSAJUsp65KsPZs/jJiBNqb21lXEWzSZEvMc5BUps1Uz00
thH8/MktfTEBEiE26ep+EF+Hp3KdgSa1sdaX0gWriGuMXQ5Hox9IkLFqHLPFNwzQ
Apxt6238tUL/avxd983CDIn94O2jOv7sQ8Hn2IapH4pcU7YRY0PpQqJHYFAfRvSr
n9+/P55SbVFe34mS/yrwOiVnwCCeAA06OJpbRQhhkgPHki+4mKWCUQIgToKu4Jso
IA6cHsAyYMmFreibkoabJslsjlnn4HaHjLKBFPT0f5zQ44+vvXXCSgabUWqDSUkz
MmCeE60bsQzc7O0HQCbKwkdDB8gGQt3RrJv+ai4iix05qZOeIidH8KEpRU6wWcqx
+74gEiqhbQH9uoxFCQthy5PzDihwTezzLFMRlCA1B7hY4ZUm4+zlQhi3aQmE9mr7
ahqC+KIApm3XVmiDywsBZQSg6jscca4E2Dsy0jh49JPK1+E7LPYjVKIqPsBHfzGF
8DEqVhWjgX0ooXb2cblfpFcsPsoC+P7SusoK0f3O/oKRHqQna4HO/lMoCg6Xknx5
+hytgJQET6fLiL48xz9zZw7LTXknBN1uSG5Q+IzkEeugFXRbiddOVZB9q3K0apdZ
qnjjqPNAv7AmZx6FOx9El1EO2Yqvyxcc71sgZBt6kNmYKmoTGwTYaOGZfw5E9mMD
kFDBPaPnBrjriFhl+KkIJscD87OOEjpvlVZdIR/Ovqn2JpxupIYM/v/7r40awMYA
OJIieiM+K27qtknouVgvD9hzrWjYXftmLDjucPkclZyMLXuzqRleIMHPIHkffQdq
z0puOBJXeR1O6gTqw9kmG4RELpjww35mirbpyhtESZUGfTY+WNy4a++keASHdut+
cK+/JsYuKZOMWdTwuEorAwFEYDc214/dKmWkcXKwtnk2Yt26O5bUqYrm62ibjgdw
QOK37cQJ9Qe5W4+pH7fekUk+3rjQvD4OoqJUN7ckEXjDpbX7M7bR3uMVY7zFKFFe
sNaLysSrDvKtxL/N0mWQ7y9vCtrtn9PyOXEisl9cJyvDf8kM7h36qVO20JiOtCUk
izF5pwnOjuOFH0Yb89KC1bffnzKL8d+LOcxPyqusHnYPmsODXziG4D7a/zWrXhyT
W5a+c735KN7xIb1z2uboq+FIgQJMQcwKeDALuQgn5vxQDB1KWVTiWVlFo5xVnr2Q
O4mYsC8gnbYb0cT91BGL6FrAcqjdZB7qmj+Rw3ULPNpzpsCW9Ijp1NSNwQ9yiVA8
/iqoy26aOr/gl2aZOSCSSR7nIBA0n257MLhz8YUJqfT4L09ZHxScFYq+Xjo/KYHQ
ON3LALXc+c5SAVkftbV6XqzSHjgcCH59422BJHt25wXRc1tcssSOHb9KCWl+HPH8
xMLvy/nA8Q1TbhW3Thd1vEQ/tcOP59ycHtGu0xdOh+ID3V7IcSzaGRkmIvr//eoy
kWqFWdL1tbLHftTxq1L8D8/Y2Ee237HlE3M+f5PoW8oretueZwrh/toYVGHWoqn8
1CXQXdkYJS3h5O2enZkbcBU08+qBQpjO4mMEnA7UQQJbIapM3CXToLQoIYzfhBM+
/hkqA5mZfMfezOpRAB6S32Qa3U+9UUc9YCR/Rt9NpoFt5sk3DTdLC4aPmlS9PbkP
aB/ZPEpENtlLm5YIeYfzOD9AU1tNg76CUwjUocXENgWHeddVArJ/N80wpcgJUzX+
1M/GlS6xTtB4pgr+4HLqzPgXrCZoTPqtStzjmU86VyZNlOZ9y6AWtcku5R2Z1kT0
VWGCE37rtS2w083a5W2RBAwIlSXoWN+s4VugHjpE75FVFz3GhEDOAzU6TFFAA2vh
GYi1N2d+Cnpvvk1hmyFBdNT+m+D04stgZLvGPRPVTgtXQ/VzWtEYoVIDOJSTHUmX
YycPdgcDoRhsQKMGlHn0zb2mKAZDafZGoPfbD3atckgKVHgsFrhB9xgZ8tN6OO3b
SQx4Efic3wOZIG1/tmdtq9haVQf9x56kyfJJq4BgKHbzBaivae8SkN2n4aEGefjW
3kiqRec2jdabskNO0tvuqSQQZdCCGqTOhSycgK5MJqFklbF/TWwXfVaeibV16Sfp
JIPv0AStmWhYyycL2FxAcgLFS8f7eIc0z+ThwI5UvQ1cZiDLgK2k+v129YMUkLiw
Th2VvTaOddYNFCfmDnEbH9f+/acXnqiPWCzPvxlf/XUgAESsn2X1FUv6sTv2tVVf
1u3ygTTMlSF5M0YvaUe5mmH7RzyFkrQulzNbUpiFkQlU7Uy78ReUTh4SlgefXR5F
r8yGBe9pRKVkGUuL9t4tau1rMEiedYOE7ZGrwekdNcmX5+4UKwhKhjxgb1nOgCdt
lfjUSR04t36yH+jJ4FtAs7mpC3zh7rWZ6sDx4QGZTIgmG2hxuxAtinyrR1lTqtBo
SGsnOppHScI//PqcdtKaQU7cPUIuDVKlEVxzhkggKVdNGuQkd6hGsoyhqrEiD+Bx
6S6xiupJdxzEQgvsLJvEApltGj0xx6Zl87e33EUNy+Aj7NEu7/nx/JdNQU7ZhupV
fREGJm4K2uMAgmQouy+Nuxs3vmoVmDGn8kwo26Ry9wxkHeXgfMJ8TFETtDwXaRbu
UPHvYMQmu8gDsl8Tm4XPHt2lMMmEYnlvJpFpiWKYTuNBl9mHKkxbeqxUanrT+9vO
j8R5WS8/W+djqG4/sLeOcUeV+LHVTEPM6QlS/l070jB7PqryybQuksrwA1ZI7GE3
G9smvcCS/zPZpafP41R0nbCopggNEThfFzYuGmrfNCS1yvzxkT3v/zAL4Sqopnli
ENiSPQmYh7kxOHrMy746Z4iFyY9JC8u79TmOoij2P+3kD0zZVueQL5bldfNESFXU
UBA4cjXhnZzcu9P3h+MsMJ468Krfqz2HL79pPyLeyiuO//RIikC6mfXD16vIhti3
ByEoZp36ZOnwwp3lqyoXRa62Z1fHXrnvko+vwaUGN/619tJrYBToifRiRA4zGzJE
gEUVOrOZfqWsDbTtS04/ZPbkzD0hRxBGr7Ks9oDhlqgkE8TCci24rIh+SCPae3bl
ThdATzEENHHijWFyn/eByswDykMnCeRfuwbLm3L7isDgOEizieaaoV7rVuks+c0q
kRrUYW7yl2U2IWBdNKNrE5N0xtnXaxfoEHGxEt7wQP8LkJSzznqkpWM5SNpSaPu1
vM2dwR+KZhZt0zEEE/AZuVzQDLLpQouHHS9pGPVopTBwkRac7L4fEGZD+/izX9Tz
be3WBOkkncA4j0vFFkFtNWUhhs8715Y0PTRUTc3CYv2b4stroG5jnh3VPvCC34/z
hhWs3fpsqmRdzxfiEJwHcCeGfLeZjHNSWx0ZPmvMN5ig1dyhOl42fIrOMMfE7k1s
HoU3z0rCQe7OflhUDJ0PhVa/srZOAcC78rN2bpw3VDT4wQ9W6A/FzmGQ+xZ5kSbL
GjqRNFO9kpgTHlzIFTZhbMHPadiwh1iU28rF5jna99Flx7bwC/tyzh5gI4zvBwrG
9uZQt14Wr/xMCNYZLmW1XNdKufBoZ7wzzS1geewLNcM57UX0MfxfdygDMfCe6Z62
5FJ3kM3GhbYl4Xh3jy9a+TtcAFKGW+ykK3cHSLg3pw05LeD/GO+vl1xN6rEE7XWK
J4UqMi+QyTGG9KSdwma05FUqhgAKuu6f6aoNoXSt9ku/GmfifOmO0cApq/m3Ciu6
lAKZUukeDMQZbz4UWBLbVyF3PWXcbNavbNrcrLd7iSiHBL9bHAm4fJ7wbPmFo8/n
8Gs/m1/+5aJWNpVTu8bPaS4RH9OIC5Q9ShsmU+i3rJUU+a/wSgwzL5a7JrH9ONxX
e6fbPRpSgGITChAOxF3ALo9d+wrLM0jlhjggXTEZfVvdhQDoFuIVyP3vpo9ADUMh
ZsXwFJYlEZc2LonHYTcHR//Tfo7jcQGXpn7kawnhw7VtZI4gXqVMIwNGGaB8adFB
+v/dh3jNyhQv62fnr2pvn9kJWHoTl7hBR0HMZ0nBvM4yDyjEFrVVIMfC+Vm6u7Pb
kizP4CUmK/nsK+zRgP/1EYQ4mNkj/Hd2FekbKye0Ubaj+sI/w7DCOFdIDEOcYDmU
KJiqi25J8ugnB/Kb3diHXmF5eX+gouKG+cd+K8cC8qA0cRGVU+g1aEf0sg0x0H3S
AoqqPot0OQ8rWN5GZ/ZMpcKvmoN8WPEiADIBt+mVAaRniz4WNPdQhKIDtkMZbk4p
RucHJq/Nm3gN5FI+a7hJu89F5tcIJXMYPlBsDqj/gEXAmPutbysy5C0B6dRypYMt
TGuFoKes03iJ4pmLJXnmfk0p3w0p+1AA2a0jNbAyRL6S30fYaG4OizslNcTp1i1W
brO9FGt4kJtgrGfRTcYUIAgXzBCrObSCUcD2/eGMZWEdJnp2XP3xbK1TIcMqdnb5
YaaXN84Fo2C55ySJmN2cmcOWRQjmM3TARuusdHFMrzcpgSNpvOwhFVjXJVMEaN3q
WWwfW0Bc3BKQTuvUWb0d2cK9MOkvGowqe7F3/rDrgOX3FKNCnKwsTvVYKatXK6da
HI6Lc3Kd1/pHlils4DWiWJdUlHl/zLn7B4IzUqymOrmvu6KVarYLxSTi4pUjiIHC
PYC79A5v8CVTvQAPCmBE1MWlrj6GCy5r655IqVebh51ZOOrG+VTDjFVDThi9tc+G
y0agUhMeqt24NYf7T4EkFJqY+yeIE/pScy1XOCIn1rG0+s8yl5sL67ZpAyHhay/K
leJLFhaWy830ln9p4niVoracNsnxiv0ahiOuCBPhDW4QlgKgV6d2wYi0o6ewHuQQ
E0z9GHw+QicMRAWexZxp72Zle4yuciir3bnNf8Y9LZ/nHiluOA3M8GTVsE/rTMM6
YzMQE4FwQUMj3mkqkvtjYJMECFbSXsP/9i3XXbGSUQINrgZIBBSaNynsb7yWphSu
OpG/r8kVj8wwccs+me/hZoT+IVisAgFruZX1TqcjAt+J2LvmkA3qkRipM/Mu/Z5u
m9XRYoT1BKiEC+xiO5t/K2EhQQKHODwnJ2oIqRjgchJ8toaBqSwWn2f9lLUczU3s
fRWWo7ttjzAq8oXo5pzH1IwcOdJAaNQdWwDSlnxdM3UjFTHAoe7TA3vodIY/IxZH
fO1o23eSBwSiFn6xDahhdUPr1Rv5vKGG3O0t9MOmAta6Pzblf8lvh4yQllHZBzs9
E7AxZ5ukmWvUdyuv5vj8jsbTkUixge4RT8hAuVlZzkcTyfo//g6/yZZd8OaW7GuB
7DUpOBZgfgKc1atWLGoDrVrBm6BJptB8+KXHboqXS/Xhdaef2gTTkS9i9ArTz+3r
RR7SixUQdhIxg4PIorheNoKgTj0MrRcamd3usqJXNY8Ml9LGJyB2MMJAa6YEzHmA
NEGALmsqysFHbhnoIGKh6rJYTkfUUXT40IO/RuLEOxBhsKERu0qU+GSxeR/GFwVz
31To8EKHWLU1IPiVccvXcVIZ7M0hu1/HgfrNLEkI2NwWR1pGPAtSy6OeOq5VEqXu
uAPSUx8T16JSCaiLJ/0iWFmHmaIKi6Mgz4Ue5eAsVKd24M1KujrFgK7AOUbbbImM
YhVpqi7DPwzTpS2OoMsgByj2ro02Lb1wxUCSW5IeVEf2zyTJPhaLP4OjNMOkOABL
D7LDyMF/km8KOTO2S7dPy9zQlgWD7kgloAQwN0r7OvatqjJRyNy4/2HGA3CRDsT0
BAhY7QtOYhmHOKAYl31XnM9kLPDIwdP+FzqG18VZkupd+Xms0ma/n1kTIi7ksvVR
YBpgimFm/ClXFGnFjjmz4e1OjlrhObFeL4hPpyh9JglEYcBe2HnHlkJfZLxh7TQU
xuVWe9iKslPn3gop5y0yhxYig68BZCSjeA+HQM/9lavFdo8QOCdhNSGqEh/dyDFS
3Avu5aC+jVUaV+ii3ux+sQCgRLPG2g3d64dMSfAgy1E7pg2qidocwbOisLadgnqv
8udxM8un3ErW/MYkVol8y4UncqI0O4yuUmtE/ch9nbVTKTC/iUerD0hOIqTlBYLX
1kjO1ZfOfHhS9INC/2ZPOSRumuP7Iip5Drsu9O6mJTqbmho5BDx4QhfbHABteVDk
gstdOQEyhiYxqOKBy5C9QCHFnaN8Kro3cRhamV4dlK8a01QLeCehD7FSFP/jLztD
N6v+k2GpeJIm1WHHzFJzeWfgWO53kfM5tIYttHQUgrm4RmjVXAVlu/0N9OX/peRX
1LDRuEcEB71hFfhGd3yWBhgzGlNi7nQrJ63u4z8GeJEQWLuWMHk6rRLgtXdRxvOT
EHxgv2iYLLa2cvtmj1CXbM0C3zLngK5GNUah1L9FhNg9Exy5lxG7Y5gSM0xLLjna
4Q0t1yrFGC3YMEz+Pk8ljSJE+rIPdbANELw8cb16UczVdigCDh8IK4jwhQ/m44uT
9FO83TbDBwrvVWCeaJaPjxhfDLKHZth8eMykM+YrJZtxY8YPQAWE1Ayz13uF6VeR
+ADReKaD3/7dRTC8Kc8DbfsVebia9AtMePg/OgJiRqkd1B16bSTtqt30u1uZ+3bS
jXyYLd3AWW6pGTkXDH1QNm6SNYEJpQhU8C5YCJEmb/xqYS+sS6fS43XZmltWq2fD
ijSMCXfBsVMe96j3JEwYCMlUxPDbsfmvDJJfiTaV1NYM6JAxRQLDrMNAgzuKN/TS
ZctQBGvHEs+l+M0gxg6Y77gW1IdPpFTMj9vvDQ9twGPjCCaUitZ9/RvzYkD1zhLx
x19ZV5Okm8R/VBH4v3DXJUUs865nqoDI7xvvcKgytGY883LAhN2ZHv5fagOiG1c/
OXb9gNPz1KhbaGwk0iRnOb8rO/IRVjs1MhtNeIoLzsELM1Axphg6OjIhHEtEHr2M
htG+1spEqCsLsvru+BiDCJZMLiC2Cj+oM78DI7tRd+NF8aWseJZqQZAFQW/xhkWk
Tm4c4UCsJKv6SSrMKBZ7Ea2ymXNymi+5xaiaako6rVoZhmg0mlbXarxznuCczN5H
gHoXOUpwroGhwWnZP87MM3vO4WmknYgF3DcvPeIrG8gbbdzAvyUyLkvTIIryx0HE
9gjGkIhtrcdPPL9brrDvcOzMw3p/Y5SxRFqnlgpuwUboQqBvM75lOOTiTIkWnPPz
mhy4gwnDLfBmTdcJIATEXUbaXTAs16OuveUwdAehPlxfZ+GjfIPEENLVLwRE6+1T
Od+5Bo6I/l4JmKp4UodUegaHaVjQJdQpDhoq+9EelrGHLg5I7FVo4v1xMnyqWGzD
5PKteI8S/SNYabTWko2PWh4hwoEW5r/kAc7gcnmknQ/ElyYCMOW6gVZIrWUJRx9A
f148KUFs2qgkZPXpmQZPDzIauA/a2xDJcVh/QKTM24JIWirODUIH6yYecwNNAnDz
FxK3rhNbIrsqaouRyDimAc497D60ywJB/Hh7UNreqb8m4azRA9XFF8KUfEU8z6wy
ipH2NfAHUioNnEGISP1oAmo3rNQK0zjdGix6J65RDcEvU7Wo8zkE47Ngp7JhYIvI
K2uNwqzxlKoxfRfpzBtJ/6/ijoxjkwunVz5w/oxvCWW20S80ZgIOsv0aig1vJboK
iiojL6fzyjYuwpC/9pUGFg766kA+p3gTDrbta30rLPOU1Qe/jtoCNDtsjzKkc057
1xpcVYEuSE1vy3HaC4alAyURiAbbdoElkpnN/vJbrEBpiG023+Rzpcr5MqY85TFN
K6XPh6yex/j0o+1s9AI9wXaDLBhfFyXrXkM0VoMXDTOBfvQyj6QCEHrzuR0JBdcI
g2+4SfvbYoXwqX3RT6b7gB2SpTP6KIJtGOp3NKVxDzu6gv+/7S0feR7heNdn6M4t
mjWx71hwhGgd3AGnV61jEPj+42vk6n0HiYRddPP/oCC5aepgYAD/ZR66MHAZpADy
mO6IoU2IcSHj8XIyrSWEYIkcPuTQH24TJvmXC6M357wyjhjiCSYvld0wLFuJ6mvX
BZ5C4KPJmLQFslFXcc/0J46XRnzdaxMA82DvBK5O7u1g884MCf1+5I7rwZLdpD0C
x/kRMSlyH/t4/mAhdVNr1M2z9XFrLUJ2EIKc88lb3yrMDFCBufHlQZUQwB/14Epb
X4qy9R8sjfZ7yAxC/gCaHovUBdG2+2RCOneOOOeCyOegojiVUkj8mF28Acdnq1/8
AUDLY9MwySP9GD/3AM9JcsSTeQIZGhuhkdxFGUBJTeRcM0g3cRZC85pLJKFU2/iP
05f7QWohv6YQOzWtdMnlZ9Hxj1CD0r96DFkd45+5Ef7V6mE1pAIC+DqTipdaIk0z
DIG2NXYJYkGhlgY0v/+yOr+2MFEVtfSV39hzgBTGabI8DHoD/8kTC08TAqOVH8Rb
n7NWeEPgmZb4rWBWIzWiytw/93uL6/EENMb6n3wWhSpTa1epDPPNORVXMYlqN8Zd
YeyyZU815HGrXTbnny0G9OhUUxA3q8izv1LaTjF92ttA9odNCnEY+lPWSm8h/2ol
jW4B854duZ6n+nj4ovE1ykAZrrAZzL/gkN2qZEOR1TC/uDQws3bE9OmQGHTUwZnx
0LSKoAbASxb0LLBTQmbdz0UutvM6lSPyQKOg5sYIBIRB1ORY6ZFbdf8MJfaDOUuv
Zo8jnS9jUGUwYbnVwBP3/NTp+tsdtj6Rvg91rYVUpcAwjZIrzKWgQcwvb6PHBGYH
hmPEdGuPLUjr6DjTt0TMqhDaoc0w/H3daEAyegOBT6DiL5OmjPzwOiclG2ZwWnyQ
uqG3m4bThXZ6dKmBe9Ar7gTAkJ+bxinQGMbK1kfuDYnZWKKTGsqaED1rwqooL1Um
Jip9pcniQPNa+9PD/kcK0OeJrxbO/r98VstT4D9e++1Z0aCnOs6UCzjMLQImrFuv
Im/9QjkHDcM6xKMOXrfb5gqUJLgaz26m1sgbktlXo4M4j0g9zqU5jaBRbQzJZow8
BPsIz/AdEz3k55bdhf3DcjEgfAAgAlDaGVSWl5NLQr+wNMzqjHUzZJQ2hJS9vYTq
P7UsWLnslLkqlreJoRQH+8xwFYhmJMJNU2TuFxODsG2v4cgGVmV6jhKIWaqUi2Pf
eG52p0lUHW9IiOMTuR6P0BKK47zM0/C1XAO/95hH0TitVBvZd53IfcWAq5vBouHc
djjfaHmH/Jvv22kQ9jcNLLPnE8uT7I4pbAW+KtsjPBWialNsITdIMVcc6CBM6zTl
w29F6Rf9WcI9017Ymg5s6fl0F9uU8pJ80HUWTWsDyQJQdKPcuIzrmn0b7JG/DsXR
yT3HYHgZy1i8SJA0W8rCsLrk5igrdzmIozwjXoIGZNjoyrh/vBbh3AugFVkX8HJ0
N8A8LwWFGTzd37BhJ94/Hk206Rd9+F+SPDUgeoxBDW8hmiBIQxkRGj5RrLUi9122
099LAOWNQcv42UE3zndsiNW8iau7hdrMZSU4Q2AuUUGXmx489oC5emoB+TehCeka
bTgZfiWk7vDw8HU1yLxilZ0Ook82yXdJslKmjk5ojZz1555Am4GDEogT6T/CX5qp
IJ3XUrRNatV5KVfsG6AkSqcu3+0LUQ/W5XbXi7fxg6wWxSV9uAXcm0C3JfpaOW/t
6xHd1lRNwdbytdiN5nmrWIaCac4DeKZLK4V4w3Sd1WI6bpBO0VA0GSX7wchf+4Qu
1WNEV3l8TwP/fZDQbkNhetfb5STU1kyMLeRbuKK7JypaUnSJVP+By3WeCA6eqGcS
4/9dckkC4Xx55pbHuLgkr5OPuWplChrE21fAxJ0K2wlRpz/0unxVxTrpMUseC64J
PUI6vTSuJu/RWTEhairraqJNL7pKpPY1Sclg6Adq+OXvmxNtFvYfTrnls0cnT8G5
mvGy90rwSua7TkG8L+5bK+XTzidu7zPi3RHV4rKaAcLfbxwURooYCEMo5xw734ua
sWVDIiQc3TGZFHHkK6ZbL/rs8ViP3XS0eMQpt5POTvxbPpkjYbSczUl+9Rd3mYJ2
5ijl4RKNT2PRbbQJGQGbjAh0fqUawg2zcdM/in9sTRXdFc0f+BUi6Usk8fAH2AMv
kqt4QuBhQ2q4C4VbrmlaQCHDQjgWr9jp3JsF9xmC+30MMcaQratitHinvcK0Dnkt
HIhmCM1fnQnV53rvpLiEu5ZEM1B5TjgZnfbCfg/kiIWZe9lWY9QI2jbnICsdc3+G
GkpD8LgenXfnlXe+4S8pSSYp8enxeMLvltleYVxsqypv/Po+tZ1ScEEz+O1ngnde
RsgxkZmq2jHMYysA4H9rUiVQxd5EgfC07a7oEOot9kD0gRLh2pWYGTwf9cBlKPfK
z+cS/1YGa+ZI2UAH4FkkDAizwuYSGr9DkzvuTLpSPzAKgogOPMh98BHS7ivVUpfB
FKmKdXehnSp5J1xV9J67cE0qBnhEGH9WH7Ps847SsoQtow2RWHBzBSd2kgDn0jaU
v520k70EJtF95KZVsRDBf0mYJy/QPf6JyNhdssyomBfgTAboaIFaao9fZeLB0prA
u40SXwoP4pa3MhDVQL6cMsQFIQQQ9yUb4JDzUCt4PdfriTzdvwXU7Gs0fAiu6l1D
asKTDTfdqCKRpNgu+KhNSX4UC56D3H3f5LrYsH/+PPDYTnAv8FomDeXlh1qHKeu0
U5VSdJ1GYGC7/NeJ7dKR9950xQe8zRXwT8Fh/7THzunSgJ5ZhHUs/05c/CPZkSGa
ELyk0qjYt02ykl+BOe6c0vrGaibcilSeVXMySqzxW2C3LoJIYxi2hN9aFt2H/qBG
QCUuJWY7EVez/iLwtcJqtCuBEUxNphnfIUH+cZ30fixSKRozsB7hqI5tH5nWMhbb
RVELc3L33yoMDKduKt7AXs6/oj7JRjuV3kE03nQfzCmQ4oiQtvRoYEYyN6yw8X2M
lMUyu995GlFVM4gdCxTJ9kzkTa53ZFJyGIOtpu6tCc8I+AiYYiHH55YMAhGQSm62
Uz5oPh1Jwqd5gvrylrH6VH7QmbIcKxZMQlk1JkOs5wfSD+mWGUSuTrtn5Ed67u69
kNXRGjoHAw2eImE/Bbo+F60PyK4s258MVP+x7kOPo3l22Yy4GbteTjgybs7tnDOD
Sar2aFG+MPnYKX/lmxTY2N4SN5vrLTxN2SE1P3AWhl/dDdFcnFbiQA8E54NfUflq
ulca3bHj49uTmm7BCzuu0np/37n175Uxzi3FLfizbVWgzylbn45QUjZ0pjZdN4ik
hWgBrdsaZqYoZ4dq3Ai3n1CLmqNoXRxn/NntcLEM/yTJe+6yZCr/vBRuWxHIQDh9
90FQfCemXaP3ZE1zIAPoTIUNrOmm7iij5vGQNUKqVspDMD5RoP88RI5dSZLmwFmB
Wk1Ow27VuHfZGPQD+Fqd9PAY21T+fCIiZTMRABWUvIfFayMi2pcMxZXaD0EE+jUP
j8JZjGNEoOwP84Epkl7+2RiuolhQm+0kYakdW3XvPpblzFkEGbAj3p24euva16N/
2YTCli9VonZrWcTiWHmLNdERT28p7SL8W640qDooPkCXUhTiSJ0du36aQi+F2UO3
ExoO5adzNbqM2IrG9Gsk6jnl+tA4ugy2XNy1k3YSKcfh63XG6fwGz3ARfGjTMSBB
g69bX/2w3dtR0WuHrGlFho9Al8lM+8/8jhaPUe8iB2S/VEKgIGAYVS6QuDplhDEm
Ywvo7nM6yv6e0OoQ0SkjAUJkX/0vzu63RfbwGWnNDazOj0xMyTFB/Uwr7MKPl0+7
x5CX7ijfDrPe5G4MBNEK8e+5wWNj+x8xWiz7dA4bnpVrHBpL/mNSSihUCHUMRiKf
/EcakzPANQC5M9xVLsJeXyeyNim9gU31sEWO2Olbzy+dbd/ckXcRPrK0U3rP2vIX
ZsX3CuO00KFG9k7GqzvGmqjM5xII1s/3kVi4MnEHTnuI4ZDvezspLWQ5FMrehrgx
xbftr4rJxsqY1LW8VF1ztNJWjZpIqHiykJcHQcg2uRj5jW8eADiy3VqBeUSUKkcu
+PAKrxQy9IT4mpf7KTfy/nkixmgTXiQfoXiyDyRsi/9n3qg+pQ9y0QbxvqoXkER5
Q0zLuAWpGRGJZmSHZg5JbjN2bhlIjfS+09K2kXpR+Am7/0RsjUOLamSQBTcOh58v
B/KjJdnEwVt/MdVZazvW+ziD3jo6E6mbESWeyqLSl6k7L8EypPwKqGkfO96jdQ0C
jULGDm7R7G/m3jPrQsf4s+818cycHh0i7mJjYqbYrlEhGvfvZF7iH0jEBpAray+5
eRCev1LYjCiyUyvOpafpZIgh91ixTbzCgnYoKSXBhDy8phFQpPVu0hJZMw5rXdQ7
0MHDH25/nSUuqANNfzGYZB7iKyrjd+ejt0zlM5JefQlyvjcOJNQ6L7nGyAnbB53F
UkFA0VFM2F8YJwiyzpXz4bo1POhyl94XpXh4nndZc5jSviezhQSd64U8KfSrFhI1
4UZUv9T5Du33GO51RjPsFTCM80IstGbVPmeJnOeE/tvglLu3OggQvy+liJgsqRhC
VSHKq66pyCFKd/dR6YndccQDHC0j/1FtNA+3twXvVzvkeQdCGe4DNxw42YdnEfdv
loyYZwSEgZlGE9An1sHTdBtVa4iIsyOxCzEIaMm1PFaSa4HhwNUUcweHeuJN1urI
5tfbgOOsgkSPcqs8ejwMqBEdyzzgxFKeqChVnd346gQW+000p7uKK+122+k+zPt4
zVt2MFH4qgyrYz3u7BwAV76Zra7PEGiceUafUogJfLbBZxytw8uyBc5fIPLo/tzb
weuGHSG4GSj3le4WM4IVcFIT3aEkSYLRqbG5zvtDRjwmZf5eCoO/qlFla+xMzW7f
4aDj0a/PDLhTzF4V3SuW7aF1y5QTCbjzOugZx37hwzbqogvJNxl7+SlOWgIMM2Dc
r8piNNyNPIWvEnFc5g8gnXPxohCGAYSfM1dg2muF1h25PObz/4BZDJTDohudieZv
iDTKInJb/238JO4O423oZz/xH1vGf/y2GYZykzgrusxfp0Vir//s3/T6HGCxABBH
o3Rplw/GmyJy8u/cx2JFRNVQwbp+XoWqvVEviZ3i8D1paR63TSRpvSd4ysKMMzXZ
cl5+G+OC/p8APP7GjiRyZfIkjD4sm3TAU6lbHAAixwEDlHVI9zZxDMU1vW/G/+tg
eJmob9GyumtiYQ0QfS3dqdwJyLfa5mr8zI0ViFCO4DIoBbDrFabjthw7IZKNUU/s
V8b9dTrEWF+wA8szbeqxWq9Rgu/KzVKPsCuw76p9dj2+iqHC0NtAttNI1qqdxMfC
UnkhRkBSgWNZUmm+jrJLzrYZOYCGL5fNIJdIXh9jLvGLon1b6F6OmnVVPXim2Q6c
TbTkB8R5GjciD3XRom0vDuCpcZM3cAwbtTg0kXteWsaDczDHSFlDY+qkgGrE/CL4
xyxHoa4l1wEt0wDAI8i0/I6fXT0NIcoo7SYzyZRY6Z4aEjKL/3lt5q15jS0mxPTW
m+WdyDdEichNoRKTdDz3t98m/b8Jbn1RRvEUJx6SVuOZbTq/KjptwCkaDlZgOsVg
tjSOpkifNtGYiqjUve5Hq3q/Q+MQnQXAf/jbgttwZ1r+7mrAGvPjRRbxuSMVDI4z
V8Zq8l5Icf50eaJaWM9rXs9uy34pXu9HIsKgfL+z1m/RK/Kkle/BT0PNhCxomrug
gMsS8BunB05k3kGuwPC5RN1WXindaSBhJ177K60HUd1nq0U7t3pCfXzEwc4jXmmR
HW/KgNfHuICA0oJC19VM2d62NoDOBGFXkkU9JqM9ZJIM+Zqe4HwFto6cCRkd6s9y
550C3kHQNy66N09IINMy5Zw5Sby3IAPI6mRMoJ8CPkG9EfEi8VBgWutT83Cgz4QQ
ZZRaIfFiwcXebR5sqbu0QXfMEnQx0tZmoXSxgV5XDWNIO5jK8L51IcX2PDGaVfcR
4sGX8isOcr3UispOe3esziwFlRtVEPvrpgpwnwKn7Bdc6O39SvOCM7fU+C5kFjSM
I7c7eebIfb5Xx1invER6Y0X9PgJIcYGGFKOjLp2NNw6OOeQHqjA+WYRaumpdeOBx
Txk57C7ZLK3UezJpry225VaiwtGfGOUq+P/wsuaYt71MfiAp5r4mBiEzW76Eg9yJ
3+50Qr3911fkAs04DIKfdnTFVuAvMAahm+ThCvKXJIMD8xx26uFEUHQzzmHVHPB1
Z6aBjhXJOXOREtf7I+I6D8XC+li1PnufqOwIKgXegNWj2/JYB/Bj5RJjnGO0MaJF
5TYajvzCSyNEiwr6t3KJVjc6oLhV2/bxcHUjhy2tRHe1eFNieGFXCo5DFmuSUNh2
U1UL9CIMS3xqm5E3v2/gQNPL4UKVVKEuKFsT3VCpQJeGgzADRFJDIZARzIvwXuFe
pbDhd3GPPC6qWd7VA5bAWW2osev7NxtzWohI0WnqhVQvNclMhx3nfFQ8CZyioJLE
dFUMYqZm+lmrcGn037h8j4IN1ABfy0Dq/3SOUMeNcSNbIwBt5XowSJQtpS/aMf2b
VCpdAmpFj005VixjfG6Qg3Sf0pYFpepw71Avg87s8npo97eSzcpqyLq9yzEciTD4
t8nagd2Nw/O/17mW6RGvXLobS9vZc11P93S/1BKZtc5oEPSj2FAReh3Wasm4MZxl
yfVwavZeblk70u7JkGrN+0gB6NpTLIEwNV/amYaNyb2G0G2Zaubjtpoc62mybBaL
fp8GMTNpJXRtb/BLHvQAYT5P1Jzc61vZoAqUsITK4fzM3yMrFalO7iNN05tnAOMX
pVpDawzV9Nw7l96xowUjaUlsGPwRjGHurMsxVfCcHgH8hHPfE1Ww/B1SdTvWXgXQ
C5P1nrvNj4UUMo5a667DZzZfc2Lr7adpA7cPDB9meN+JMsKKW4p8v8QcrYt3rIqy
/Im3jVjUXvIZz8HUFFeSuFaSNG/sT1Fw68PdeOpMEiY9ecF1eG2uDEl4R5KRkyvI
G3y+8cNIjGpyksmCriLXnP8hnPxJ8iVVzTj+kq6BWfFGGBX8zQlFK7a758OEuMkm
5aF2oG5XIgyci+hO6JapfHedyFzmk/5tWkYgp6uDy6+fedZ8n2JLxVaQEy/4tiCU
5D/lniG4XLZtWsdH2QES/Z7xte0SvTpyfFqKXwwqbhY+BhVaeqmKLK042Y5VaIQj
0KuufwHa2eApDvZRitvTzbwIQsZSOTbTT2H/EQWBxJd0OckBsw0kL/C5Sfs8aFMJ
9JMolqjPMkHIWsf1eJ5ebCpeD5CqRTZ7cDn2Jz2CDt7jTElGpdQ3Sajc4EqXyXnQ
xGx7F62ZbuCgw0Vzcyg7Hb4wLJqlwvuV8x8Lp1UL/dpLo9sVT4we/dG8Vp/eQ8p0
PWmAFByfCMFk7sjez5sfCyJMR+AwrMvEHlYIB2OVWuyP+2Z8njgttIYyiqZACJ4z
dzNDbEKNmbTxOcvjTP7CMYotjmKRg3nV8uHm9+gE4J6CHYjT4dxrs9/ytKxEGEfn
jnw25xTjv1zmFLgqyzwL+AlrEPTNinAdCoCIcLjABkgl/5NN+mGDe/H3tQlWPTrA
wf6zp8jq57kobLBBKzyrtZvjsh5PiFlDbpugfieI/p+bT8Zqy4a4zDUIq9wQ6RPn
Mmb+x+Cq6VRbIJwWycjkGXzzyfclFhecXHciGz1BG2ofNrZOorGzLA0QgWcXCDpC
`protect end_protected
