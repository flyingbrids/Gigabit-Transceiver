`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ezkhRqUv/EvksAAYvx0y3dbyRews5unzSh6JLwb2UXALf2j5E/kTGZmPEs6jLjZg
ZkKFHRLMByI+DcWr8uqMnGiTIogq8TAzkukwd7Ebxz9hvs9weqa6ZVw1POSVb1GQ
TVj9Py8e8JRibqoyY4w7uArIvhzMK7rJWZP3z/XV/hmN4yup9ZN1m1N89MVPbv9n
xlI4bthZejcTfDu2q97H8KIPVtoV+RhO9vX/upoXkBA/5wtxNngwQkbN9KkOMnPM
L5gmyF3R8n5jTUOdsDmVCbjH2B//yA8aAVjcfVvMLbyVVaKvCBdhfeOQkfMUHE4g
wo4Zs088Ngj1ak7dMSOxkA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
e7yz7YIyBCsJAm3/cvLdbW498HHhu89TeVP6gi3oLMNwP1AtcbkOf2xvd+SHjaxQ
gDFsL1RAfJP37bHjjVRFsv/prporjkSNdxScRdP3XEDRc15VZ4TyU/KjTypwlBaK
aXkLZdevrS2IVgxhucP09veH/bG7k/Jl6IkF7TQmllI=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8032 )
`protect data_block
AMM7NO7zbZSfCLvPOYpjbtPQtFw2ug2AzLjhMto6K+vW9bZ6a+9WSBVGCf9Bf6Sg
Y9niPs41dAJcKmebpWeDvohWrJRaeJLBk9qiDXrDsnCEtAcev5U6tuvgBm/BbuqP
hoSjFhbEx1CVTmKRGBHm7/0A1zA8GvYecKpCAet4tH+3lCvgvQHGQAe6lgXf+cfG
3p5Bk0PrhIiKWWDRTIwqpeYCan4Wa1YT0jxcxSZjgu/2JOAJCAMP/j8Sj+A4lr+F
akEcLXFR2wUuu8I2YCJQ2vf80jc3QSVl348djyF68XByHHjzYsfWd0iyGITtKx5d
g8ZzjvFPZnaz1n9M0vC1nNxNjfNm6r4sXk+7K0X3AqNQG1EGfajwUAOlQ5nEUlRp
u4UA2uhINNtGzptsoJfh6bUUjs782BZz6Ho7Sbg9pJi3LM68R8FW2jTry2Zkz6Yt
rVrhBQ6Oudq/JIJBSVLafIxlUrbVWCdz6TWjKmyQwIcmwXNGa1uPZsLFd+I5cg2I
stJXq2JWtVTd0RV8IJOvjN9EBohnL7NoiMkS3scBrcBlJF1WW3y1tSnjMXo1pfwk
rHmqKQV07ApMWZ9DIbRLrsqbnWiYg1vSUf1B0v7vZFteO1rdTZv38CyRP5k3n+ZR
tOLmaWDBP6obZCSpc2RxFPealBpFq0WQKmn/47byW1gO0tdc5tvHX9ZoaDZlzxVt
hM24FFptCyUvS9QV/qzFSulGjyO9qvMJtizVyg++3TNMNwVaQi+ShhTSdKkuzvm7
+PhPLKudcGZEY2gAgzYe+ZbBTIXQaAZDP0vNbnYvQ3DwliGxjG80VSsTRWk8TLqs
42fU9JXxVeqSedIZTo6syIBI4OnWmrn9hhRaK2AZLshIwgJZy2L9W1aGJH1tRvfm
gMn3vzKPQEnJbZlQKqyyR2a3LSKB8AAUkKfCNILeSWvD7ymlsTCrjh+436RLCoME
SmWuChlfaTc6wm9dZEKImA+OqZdqcaGmzDfp63nO1gDMSljuWqE/XIH6mwVxQYpO
T2brJywnnWKlEuNMJwOXhyXxuYvvskXZlY9W0wCer6gZoR1QpPFOGpfSaIukNiAe
6P/uAHmfqCFg2v3xDp4HTtWD81bfPwNvbRUtoLoQWbkl7I3mZ/ilgDbFSnIHDXoU
ih4F8eDDHXnbed01CWBxd1dJg1SCp9hEln6PrHFxtb83OpNmD3oWRODYfw2O4a1r
MBI/lAwEXKG8RGeYDEmMjjVDoieszGFRXjGdeL/Q86qiN1PqS8Z7k0ctAO05d9LB
F3mnzmOkHzeaZEvPl0DF1ejaPDLjOmqtfPEJN8KxZx62DBs43ecsY55Htu6aQbCT
zOV0DEQQkIreKfC7pn4W+3f7XHrDFwMB2B6FZSYJSJkbC/Z5nvzJg8u8vS35VrAw
vprboHcZU0/KxosFIVj9F6d9yaZGwp5R4pSoexG9Fd6CtAosWPEjFnTCIxXNifsX
8Mi0M1T5y9UdhY0v0cwkZrxZyQ7IAgaGJSe0ov+BxSZY+5oZgMp6qETQBFt2j3an
gpIaaN/jmI4qwbpYC1EMyVCW7wu5i6PrIIJ2r3fxvehF7k5apmfF4PkpTMfw/IUh
JiPwtQFNpxN1eIF/Nsau0Tdj78VSt8HkOkybFhx3Z3eZFTB8U+vwY/Y7X/x1tfzo
FDsyRUR3rlm/RiOzBTZDQlXw/qupNnZi1PRuOS/KTOcyPhvJ+B6MqtQ1FlOipPRm
8MD4s/qq4TIz+TJlz5rFK60u27LOGHg3w+UifTJVsK9XI2BooIxG1RL46Yq0Gcld
apLq3hImezti3pqDPj7tMZJNYFlI3NypMPomGYn4XSsbfNbpnjX/e09icZXFST6y
NHqRsh8dECIeoyUg6ySpHs+vzEuChGRsqzeAjM93ih+E2NYou4ef9Tuy3Xzv5g4W
8HlaQiL+ml0zTRrLI3F5YMxIF2aqMJjc1eOvWxMh5zvoOOWi9fbmbJ4XBqxARlMV
UIIeTQzVAGkIUo0EVWTCgwhf/fYWpTJSw1hD/B2pz+RLZmFt0uDDEduCEdra1mpS
af+vm+f/3lOFND1/jlmNAOOeD/nLzLRiQ/G8ZHIcAFLIffGzjPZeuetCvLTlkdlX
d0PH40MpJNkfjsCm7hYnydJyUSMfgxk5swKkBWuzmvmV7ZvnzxbLi0oMA/WlNXgV
vNVtsVQ7KcsABUNC/VW9SDcj3dtp1pt8IqurGtA7JLEy7qPM8UkiTvX1yj8Ltyh/
XoqnFos2G6iv1EDK1mrtQZO5JGAZAE4ylHstYnttGtRlSuzKVT1U7mQqwNE8d9mL
/8SR9b5K2rVvUmPz2oIe0B1wnUgHRR4vk2laYRBz3yuO2a/Ev+plJlAFQ92C1JrD
lSi/1M/WO1fdRR3VgQb812BCMwz2kKZ6QbZEYEmyXdiHHogIWGvWoSliJgy4CNzK
HqoRbEeKCRyRjednsWVHrIl7zKAbHs80JJTWUoi9JCjZClu3i8ApCEK+KnpMCcCB
PS8dedRz2TmlfthIh7OD+LQKTD3dGK8qo/o22/8Gp2z9qbDpCtxJTg/yuwsKnPWX
2YjEDnA9gxSECGqxn4klQHK+CZugwVD9n7AVGT9k7aaECAyKdJEHP9OYPAsfE9eL
ikom0SjA+oqyGtyCtPYsScwD5cQuAf4E7BG4Zl3I8fFSsjrpz0gKP83GyMRgQxq7
ah7KGWq5T+wF7u2gUhMMiYq8OJ+SXBsz/ZvGn+eFInwp65MK/L/Vg0BhbbCvDrXl
xV0yPtaXtaYrKqe1eXlFQFwzP+mbaq6id6Rk42Vyr2UYANS7AvwlOkGaRJybvurn
SZxHAoo+QXloz4xi4YEXqPKqh8UtUZbqgS41H9V2HO5Mzq/FGwmZP1tO0mvfPeSY
E3yycqq51qQ1tmgAHLQrDX+PTPnGA5hgb5t1DtfF00Uq/m3Lh2mWHGbavzycFd3i
m+KoB0cXsgNzhQZBLncrkIv5LiQxlgQ7YciTLf+FsxdK7bySJiDIeqUkw2iXDAZR
qJQYAnp94uEBmYH/Vu1v4GebKK1RgF4Q3BW/c8ccCFRRWhrxdkHFld1xZAvVRVrj
jiFr17JWj2av2dRj7FY21e7r3Wve9EzHE2MH67PAXwUXoXf4uWa6nAnOe8AIFBwg
z/grb5NVZPhh8RIT8IjJ4Twje6li2CzyZHqTQ0w6qZ/g/xzgHSVEJWT5RyGLDhdj
7SGE6BW6iIYfP/sa6O49E+oebm9ZcfV19RE3Ac+K/YCOGaGrkSzr187MB4tRk51k
olYekO65ABhqVxhGxuWdyKXsYc7viLICl1tkFyI9xVwb5cDUChSU3RR1jI9YzSoN
b/wA0CePJnZHk4CjjWQrPHPcdRrbBvbbxLLvypuCbAhsCh/GROavSoideGtG4j72
ygFOz+qW4S7Wr48ULsW2t7xhbmoONczmskkb8xOdXyErxLRZ3X8xtj4bbVrwSOdT
2LQaYKGWGA69C9LaTusrXvaff+infaISTWsgfjbJ1w817iqDZLpnw19/1XMUMfcA
uMwYhiTr4AlUid3BNfYC5Fm/Jey3/p3N52i8DuFeb1gM3LTUhoygJPvgBhP3Apg8
BvvYKZCWAdLYKrnzv0fp38a6mgHHE0e6FIN/1GV1+3jJUlWPCVCYFl0PdaoyZrp6
YVgpsEx/77XVVi8FKOpnB3P+Cl28xSZgubIfdAhL6xLAmB805w118LRHoTAJKEqz
yghclsQmVxfI+EedE7e83xlHhXubKXxHB9nua/QLIdt+aiiA4HSP4evBJ2RojugZ
QLs3AYAheF/niWzZf7GPfKjsG5hnmKHevmN+GboSVGdw1AncZbXr628IVfciMgwF
qJ77lz9XQ8xGwsB7YzLNwauO86wx+bpa/cBd76Vbm1rcQeqJnt7aPcr9mh5d5R3h
vYl2+1ivHTRjEDA7/h41lMyA3psbQlpUboHh9RppoDKtFvp/iNbILWPaEnzAxLag
2CpXVZ8wf9Htxcnon03WeMQjn34DOwHY1NIMp0Xil2O5zUPgF12POkvs/DEAcrZL
MenL19tYAfTH9kzoEp+5QCapigSVdtLjmb7AFRTEyBKNLu+GbrWy4vTSu2iYAj+f
J3WUVYfGfEBGze23J/Zv7Ss4kJSzjx10Om/2g7SLDJJm3uZQsPEwtw0a7eKaXkh8
Zxrs/BdcCsd22hTKCx3R7VsMlR5NQ/vn6c/I8WBfNMjW9e5UfF8E0yeFQtwoDRr8
D9EjS5u9Trdz8qE4aO6ShN3ME6Ery0ZCyOi5UGzJ3a0EikhfchC8lBWPFbPh2yhp
k3mXw49Jd7y4owQ+F0rP3O3fJ8EngHKgY/EBPDcvo9YuiSfVDxhhFxqGvV6bpBqQ
Q1/sFeQR6ck5fl+wdoGy3T4cYBG7TT50Zj7bOMH2bX4dtKdrZ+FXkJ0jyeqbOGRG
FH1JrV79dFs8v5YkAqj2uzcq8rB1uuJO2VSv0LHHzAWqJFDZGvl7i8RzTB25oFih
AfXINxRAdP/UiL93UAaRFFPlv67Bxza47KvC0B1W2uZSZ72p4ss+7fWjaTjjOJtg
eY7kQleMCb97ZiRJO6T8mwKiGamu6L5FoCj8tbbRs4gvosa0nLJsJCnxdl6Oa8wu
HI/Se6Uy7d29zX4Vzz5dJoXrxaCv9Qa/LCt8E9yol9BxPUMWTMLgME0NKrVDZdvB
yetpkCYWw1k7PDlL+hJs5Tx5YPrTOTVWH14n/NYk8jC/nkQ+BusCOb1NjiRkSdmJ
EgLaBQLnfF58gpjFhidSJK7AQVdKknnwD1IHggjbp7HTtI5NAzPN14ydL7PEpAo7
bUq4vDeU78hNrvw6gcyAyVtkMEyu7XswDyBjGY/PeVKnnCPAvvzlHrPZtJat0mlc
7sRlk1HZi+Hs7zeIvhrpnaWolJUnk+ogY1n4kAO0oWnoYRBgit8OROK50Mi1AkLo
YLarOT3TC20CZAzka62BWeeDEzcHlBUlvW94IAkUzvhP43S3CqfQp2pYc2LSxBHW
vpj82AcMlzoaMi8Y1+3b4WfK64WMwv3nAfYtkcB04zh8ba1omYcP2UQE69dXierm
5sszecj7Eq/HgR8/+/dOXmtgr4OSG4bH5xcYgvYspL9UAWHTVvG8PKALcN5IXGZh
dnr1abnOHewCA6sk5Y4shQTiEBRx2fiidY6za7e92oPDnQUXpu2e9Xsi8V8atmEj
GBzae3GoXHED91aEeh4qLf66aOZ2gzqiFXfOT1NntKVie2K4T6nh1uP6TpGjNz+C
HdM/fyJUVNvEaYvcGGhtUz3o+zRxEcpGqt69bgbAQlOqSmHjgBqxKlOVYYG47UmR
OqSCMcg2lu2DIBLuFxCeuCdBoAM/vbIZebMti9VNlogRpIh2nF03RXFUIthCv5RS
8h5dfCMZNr2xw0EP+u4IiL16eT5AUx+SuDXNFcLuWq1J6+jN2O23LHBdPOzvpyPi
cxlmittH+bFGE4tdeNy7n/YYtf7gFmUNUI8vg/XkRabPm8ChWkKuSdIa8KVdop5O
Muqd+cP5DMX+mSIm0Jx7AMK4AUD65Zh6tEuy+DYUOxSmVzWzVu0EcjLJ8oV1iWuj
8pwDMlxDjsa8VbHq1ApSw32LU+eS+YO9oBMCzzM5MUd1igtKTTtGkjKrCkW8Tz8a
DKIFRNcFsXGEGhNcm3lRw11TbW12I9qq7cxMRUhQjL+HBJ9tZpTMY28ZZLNd8szV
/HIpDn9oxQW/J0mb3nfXP8IPb5gznwkr9x90KnS6ZRj5SfqSzb2+zD90smpdO3wV
+2MwJJlAZ7eTrm+hHRrOXDzrTWyGmvYsW1NK7VHwa+qcUCBmgL/q7vnViLAN9a2e
YDFpMAnhTNzSll5+WkUhjiU/NdB61aIk5xk48BuH+1EwEPUm5TMMSeorlP6gPprW
BgsY5uZ1Dnt8ogRP/pKClvFPBxByV7M9kWrp+JM8fPOPNCs22C8vcXJhittR5cBP
pLnetAXaKNp+FuL7iWqlxo2cKjLumHRZ4tKurGnO63VuT+H9WvgQbFA4Te83t+Sg
S/TwUef8gmHDiQTpmql02PdhecHurEWhG4BpUz3TqvPSWjGgc0oilW3cYVzpI7xT
7ffKi1xe/5G62q2OH0PL9WCMRfOM8tSyG6lfQszgpRwxyQrRdv6zddcldGfPTAx2
mvAj8nEHVtop8gNhvURqepMcsOmPjALGahcx6jVQ5cfenCSVQqP+Exqk/28ujA5J
CS9Qzh5IACTPt7djzlPy115YXGAlVfIzdrPahWpsbhTwIhFakVOVSc+WQDEU7LWB
3EdIjRvNOjHtB1VQWs/FKZb640D36WKl/rKrQ6/Xhi1en46JJ5cAJImLv79lNj+n
KAD9nA0V6k4IYLsY5sN5b5hL1E/lKcoPRuwFlagU7jfyOMcn0WqTUrkrTqYm+xqC
rrBspbgo2iNx/Ds+X6f4oMcmcFzMnxwxG7xnal+4FJmLpQy0gnhHQNa3fSbCHCPd
yIWyEXMbwOWimZ2F7IjKE13VsiPun6/j6faHnd63/AuANSxUorkPVro6wU01PvN5
1ibFEg8oZt8EognYmDPsRCanraPLeSgCUlZtZS7E4xWqkkPZQG346ktwavzLAu6u
cSiM0EKmufiSCjdwXC0tRzBGGUow0Lzs+b/0YaCg0vHxQkWqcy+f9xolIuaorJXv
rSlsXxJxUsjb/tj3zBPqjEImEUx7xPJaQuarto0cKXKN6SkC8V6ZR8LUDwKBXngy
cDC82SZFaUcEEJUHshiQ3IWL8tQ9GcB+3L7AoTLhE57fzxfo43yqDCFSd22YtMAp
KWzWurEhkeCkOlUg3jJBHtTHbGh9rxU2fJFsFB5tVwe+eBO1cxxyYT5CjsBnafyi
VaG8qDrK5wB2kynb6n2D4WJBytIiKtFORavIPvAZpRnQtxepM0ZnY5e3bJyoQf+0
nqVXdSabgz/ePsj7QG+T9Qhhh0x181qN606li9ojF1GCKp7xRuVazWI1bLyRjOhq
KIhYaaST+Y6fmuPuCBMmIIzt26+kXKQEzl6Z3OyJmSRlDatLL45EMNyIEDPf7c3r
Fgd9tjm3y0gLcTHSUPd5m/jrFTBBcx9mEfPMXu6LuIzc7AFwNzPplnvH7ye8aJMs
srC7K5TOFm0DCm7RV5qOZimsc5n1MRijKF7gwqF9TVdEIhbdrT0hzcE/bWXwskGx
iax2iCBv6w4jA4m+ck+o55VWqMF0azqKBrNWYGxmIRSMSNNGjqb34r5WRYx1brea
UNQqOPFwFR/2sxh3gBnCnCTy94xc5nB1oL1/5X9cScyTb8TgMBgGwFnf5p4chxQi
NTSiLgnM9KLfKNvDekTtpBO7JXqxsl1qQXunXITS8A4O/YAMZEAU6grw+uU1q5yB
pfVSN4wUSRqiZ84Q4TvXIaj+Fgvsv3lLC+NC6LAMJ5xK1e3jFo/mMWwokdc8XMFA
oaDSeNurRUtCQeTqTTuRiv4kb9XxiHtVivhdLrPR7UINGd5KhS6O7PDcWYtpHgwP
0xeXY1/IT4y7eEv02RcXz2EwNcOIP1d+keKm3zP9QNZOOMNIv7Eny8SdAdvKcDIB
uHiTxER7Er1V+ZFpr1yi7HZFC0UvEeBJB601ZCpqsxDTpco0tuTyPdvNNIdnwoDE
0lwfQc6j5quHq5Mi2qFAr5O1v1SuVrpYsSEp0rXjFdyCQTD7PSKVTf/UR2NVOWY7
oJDGqN3gItLuvQZnmdRDkF8gHCW1fljxjSc+ajyge9UkCRbAU6ZTBEJUH5tRhQXf
pZwlynqLid4JusDPNsbDdx2oNnMxQHWdZx/UWMuMU0FuQK3yatcB/P6IxVmgPBt4
ckICwzUVBL/m73LHILw1k4im/GnEXrgNrUVnF7/KIHYYJa+Vg0nZwHHZaUQxRg1F
DBRSYIMa8FdO0AnTd2GNKmG4/S0qBBUtb0E8H22KJYji08R6MmYMQgSftJeyEML3
eRwy6FGUne/CHaObNsUn8sf04zxhbO5ZLcqgWkUuuKrVlQgrnFlm9+U5AZ635cy1
cRKL9p3vglKNQyAIS4Zsr28I847+U02NLb67NU3c82P/e/oWKoQEqwaSQMloc/QL
O+uowPdbyU46EC9UZpaFPc0SjLGlRKmQtb8paYThWNIVfa17qBQcpNyvvNatEWfZ
W0FsLBSSjTLFNvbnkSEKz1nqKArKpJNKSe8hAOgjdgz9Hrw7kGxuK2NTkF+TO3Zf
SOvgp7RNjMWuIJQg5tXo8vyuri3Vjj19Rv7vZkt+oaiLCy9vqfhybkyCG8tleo/P
Ix5B2YnjJ0eux38HsSiv8TEs38A6WkXWki/s63ze/ehBzejizBZaKq95oXr82yFV
SigpIxce0nYDa5yL1C87MfTj8iazqO1Me0COQFkE5O2Jx32Q4xV2m1QqBwGcWHio
hbJs96MTl1cZg1jqcrwVL9dTxRH5rg0k9J2JRiFPKb2EWUmMyNu2cergOcU6t7Jr
ZNRpi+gkC30yEU4BN8PBZep5WJSAonFUYhSVs7913PqRL7ix2z7WFNHgm9Ke9Srr
CR0ytUhNJtu6C+b3XNbkCEqAobv8cTMKQPhdqhxHJd2IYNRFHg9UCVGfdIp1qEzn
O0uAhLySyohLvT1XDFuKjLJnMEQmE1v08yvKtzS9tu2Mz+cK1zFK67ArZ58oOspG
pqnms8wr+2Sxjb4aOOfbLcKIL6SWafMk+mZ4VFZ3aCVQPNyThEokO3LqHFsnX8IS
C3kJcRTSZl+kIcQiiRySUSnjn2N158gaTTJFUtbrQLQ6irIzz+GtotRrSUJG6pOn
CPpJipr5NAzBLfl6pYrLuYfmTfxvr4CKTL8NcFVUmDWg9SfGbeEIWCdH3+AtaAuE
KfG7QvP1HZzwCD09sTd2KyfeGOyFTHH/ie5Ju45gWWieTtwwIRHVMyj2k24dNW6g
88TzcPAxTeeD1BSITicp3NMha8CNMuy187oPyWB1G6p84uyjWV5txHJwzQZtWd5y
qO8tMi7thBLbWOqcy/o9ItEuw25ZtbV7ZLBEVnRCnpNVLiSVMscy+mEy+5nOqFP6
JCF2YHgjtkcNJ6/LGuOsnSQKgZSsk+CPf2q/18wpn1oEGItHMoAKwYxUu4GvHqG6
zIlFJxL+my50JOyJIGZCwzeoVpcRBJjNqXvfdNmamLvOoWZgVmtz78qtER56IjUY
HrWepjfOjI7u32UtxM4yhakZxC7fFqG8oBQWNHaqpR1Ues3w7ZJR2zUkeyECmmPs
mQGzOXuu2Y6HxYH9abXLLUGyk0hrGaTR6s6Ync7320zRSkH3CiSfkYD82djPbo0w
lcnYrTDylcDaY9yf1CY5WhzQSkJBZVgIMpLbCvtvbITxFkrsBpOWxzRNRhCp52RB
ZndjUs9RSjB91Vy9XxQvPKyNznNzAo7KVvF+MgEvIXA2sHzEbyjqTCJ4uxXt6+AN
1BV/R9d7rrVuT/G0wcFv2Jsixsc4Zb89iWKEy3oonfw54e7GwjNKPHS+trXJGTEf
hKPdIMxYpIekYxWRq31xQW/v+Vngax5vtxPPtoyFduzpX+v0SB27RBLq9fW3CIl1
ru6wm6V5UkB92WfEtr/RYHORoM+ZIi7RShn9pWMrtGyNgQyFPyD6pZ4tDW/0Z960
DDRH5p2/XZJyz/HvCBWCo3Wrwd9khaYNq2Y+yVZr5ul82LZK/f8D2aA+Cpk7PXVJ
vLpGzDMn2y/3QMMzCsUqXugSe7UEnIU6F+lRMdxsNSAfxC/zjXtSKXSvK354O38t
5be+AyzvvboyQtP/NL11HeWhlRmlPoQseNyR9xqYw6xdD5YyNaNRHi4R3qqcstvz
4kv9J6zuNKSRQmujrtXM9BBjT8pjfOKaCNcyOUqgKT1mO2qqB8VHV2Ckxu2CpI4G
/Kz21Hf6ZUiBXQc3A6d5tzAmVPnMoOYlgvWh7jssSkyr4SP8k6tGueELmxN3sjo4
EgPsTOtRM0aCF5MaNUucgPUI7WA2zLHGW/8kN1PoRo5bzbMpws0fjUDSqx41+2ep
JGSun5qT+pxraGP1dbdDMW6PgfMIbaHuuugCkxnAUIRQmgtyUPK54qvQVdgmkGWy
lrJAdkAW65ClnuCp9ZxjepZ191cBCXlRLAYGy3KJzCc9ixCQV/V2UXlBHjtMYg0v
V2H2DAcJx+R2/96GmjcXbR96bNKdM9RbLyXw1EkLegy7S5feIsnkhWLV9g95R+Y8
t6Nfasiut9Gh5O7At2ere9vcRJIeyrrKdSAaAlWDnr/4duNGsoKkQb2IYiOSxZoU
x84B4aqwwq/LmG7qHtTfjaTDvWxvVeU8+vjEBrMUeAl+PaL1c0WRTBeO5NVnHDfY
X/yukvTb3LnI0fONtm9qUOhqQ9lm1qVpXhKOckQzGgP+58WUoM0aLw3eCtSXxNbQ
+EdezldiuJ78nyYx98F0BXQ5srhmD4pI74FFQOOUB4NeUWgGMCUs4u43jNvg2zgM
/aappxSI9niW76rwoVc6gRU95oWZg0hb6eCIoerN5DYrNf9OINpUVei2JrKcj04i
e0NLX6p7tYQM/UOGvWyXJwGjyq8rELO71hSO9e+7RmJ/jG1QGnVqN6GHi2BZ4sCk
/Vx2TIlI1Nm0ia/51nslFHXBRXoNNQ/W1qlrODJ6mEqqxy+6sI39VZ99g80LhHgi
esGJdlcYQdLeaoRbiYwutF5rJigkJ5wwfOovNXqe6krsvdol48Pvl1gZOJQIqPMX
NS+TDFPvz1UJzG8FQLFs4Q==
`protect end_protected
