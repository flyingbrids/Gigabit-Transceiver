`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
qx4EkfcqYk6ujpoiOeSvEqYCiY9nkSWTNlUHrim2rNhHi8ZZcAK+zKEHwm/bfXU7
hpwwcQSpZYZbUM3U9+6NFUcOfvQG2M43mOfhX2xfE/gg9I7TzYr3ZkLB87Sbszng
n8fcpaOYPzrMoaEMXyphPzlpfmJfuVRKT/ZYgN7TK1gkNU+QAgeRSfs5kU3XvEIo
n/hfeu8cq6g2gB8Lvog6gG5Q2o7p/5rVfReRUNVqgS1Ys8OZtzkVG2xZu8sl43hW
dwwdA3nZEkC6WZkrVIzFlZwA1RdkFb0YdkKfec/3rAcUJRY+3th5QYGnffvzUi1S
Imbv6+3R+G4qHMt9N7xRUg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nZ2xlbnfr60YUOm7yJhcH6KVax3CvLnNCXZv8WGALJhHfDteLyviojc8fLQnhjab
Rso4OLz4gpRpHc8AO57i+ox0eiRW7UcXrkkYab8AI/XC07YrdWJyADJ6xngqVcRX
MCfF5CuHiT/ytWVsfdcoTH9cyLGmXMt6j1xYgunAFQ4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 116160 )
`protect data_block
fjv+prfXglc/yoLXhXnCDAgIRAWEAU8VTTNypX4RHtl0/ogME9pNfo5lRNrLXGpi
EAVoSGwFoCiWpAywbpJ5j9hcCcpXMb3dFpQ1NYjPZNEfdkYT+LmjXA8IIEf8u5eZ
uWxl3TAdaKxQI2zLiodrrJpfuKEAKmZTHWA2l3MG5zIZ7q2mLlvC89/pcVMcYZY9
u4Ldu0fSWYUPe6MLfJTMsy7YGuE9HMEU6j9gmnSLdJ2lXU0slrC+5lM/dMBVgtsU
tet3S6jqfrLjS/fMa30/2sN+jVQr/eY1Sme+phlX0gNL2PVhq3t0TGw6RwbxSTbV
KxrI5zpCbYg8L9EAlLyrHbgA600oJcPJifSQZTCcxfh6VpW+5T8exwlJQnoqBixv
22v+YzIMD0SDMYFIgmME4cCAhaWJcgtjUnkqPTJNfmiX0pbd6ri/y7O0txUQviNe
f5YUlcDR0QcEBX1bmB5i/WWHPxdT5nHsgZFcurLr5NQDwn+oWj6vLI3mMI1K3TOx
P5Y0NkVwxROwqWAhCq/IbnwZjs6LG5xMkmeYTtU+e36ft5cImqn+9meJUU/9F2Y2
Uqr8PEfOytTJl54xUwS8cBbjgdj1mG7wW4Ij1SHZhdl1nTUp2VsvY/tPKkMF/9t6
2EommF7MuGM4hnxulTxtsfrx63O/dBF4QxL65QbF4+tXnPbnJYI1kea/BsY32kHS
wLFf9fUBeIk9TD+TRWvV2hgbvk9vkzLY6s3UltmZ4mKRSghV7yZwD/xdMhn+na6z
72Z+TJ16lIxasmro5Jph1BZdqpN6HdF9ch8u4tSMO53Da/pMeH7LZSTTPhD4745z
/BSrnMlHbtPXCy5dUVJ7YEdbOVR62uuA27wvRkajNScnXDlYU+phizdTUR3Uicgb
Y43JNJd7vkZO7nkzkBoug38Reu+H8bgY+OLjw/JDkbo6f723a9/uZ6dcajpSzafX
wuGj/rGfXs7E8dtAJ6vnMZDCPtwXmRDOzybtGC4W86RZqYilel1R0EaTYNF39Zh6
y9bbStv9hVCx3nE99zXJe3W9UR7cUCd0iq/AkAUCM90XOGhk7+KA1Ov2DZKrtb99
pcHV8UKp6krK7tfRcev23OS2m6NSgsy+u/P4E1MnvQJHr46LWp0m3JMDgsFA9GQ+
WBYEmHFZ1tCGpdGZ5Y5YoLeZ1xUXaDiqahiXtegaVbZQsuS8J7gq5xvsPd0x7+UN
0+NSdFm0RYl/EgPfzg85sb5sAq1XGrS175F/gBY77q9K7Ygy5RS65b6iMGtraOpN
p4nhZeAHavdk0Z00ssn45gSEtVdBM/c5pXjbLb9XpJ61verNIzUPETeSPKPjebYm
8gOFnSzmZegzgwxbb3C3+SAI/6wwyhUGdD8SNKsbvOkA9ftHLv7kv+tr1IYqBjOR
KryDboenBvX1OTvluZ989oaJISw0miMVGludZsemwgA4kwxTD+FNdCCIyuYPCAHx
kYNy46WA4fS/4lZZ9wdOcL3sTKUBIaTm0CQ+yjJb/tcaHsn2JJhoyDNOdHQBEHPj
+nXAmE4YGFkINilGuQBBpVtSzx69cTIemMoWktRhq9LYuLdDMQmTbLvxanLinDKk
XxPDFOuJlDV3zpzcjqPQPBsg4b4SZ+/JJZDp4PkjofXxkHcVOOUbRA3/pRnrnPf2
ip47RTO769ndPcbr6yI9yUVr7kR/NUxN8p/Pco6inx4KS8FcCP4TpkVG50N02Clz
4mvcurwQ6rpjNOcAGCh/qO0HT+NJM+FaPhh2IcPB7qs72nhaKspYj0RlPIG9Nofm
IYWjgmXoj3/B8yJgLEWcfq9kMuf0bjeOOgXA+SsI9ymw7WW6XeGFuUkU2OkgS9IG
TNq73u/1OMA0l9z0il+Y67BKYgWmUySp1bk5z15LiNDBnFBwXg7bJnCzWGccdUpd
gpwRmcHjGtxadLf9FzqXrfcR7pD7w1ngoQvPJkURtmkjw8GCFAHXhex+Rb+EEUTM
fAA89DS9mLKkTdzpVvt5usGp4g+5Z+exwso/2v/m4MQfULPGZKw05j/WjBl1vzQE
PtAAoSLxzW9Gf3zGO1Q/p3JWl3N6+j40CjdrqnA5wIW5G61JcL55QL21/PeCk8NC
RdyzEfOreR/ryaMsEJPBog1ZjJnrYCIuM7I/2Z1HGbS37nQ2jKzwheVDMA6xg253
wxhO071pEyOpHUIUGLD4p9rWt6tJbXtoyA4imv7jPbDb4hmbVCOumnNQmwiMpCqs
mgpOW4EyC7OXZ8Lz9/Nei5XOJ7+Cv4aguYDrHLxzWJrzpsfdI9eX4C5zlYwbnuay
hQNe0VRPK2arPM/iPvJBdxQnPaoFpUidYUAJ8i68Z3SYTfPSKii6K6HxpkwikwrU
rf81PjFka2kmWlDoCgva8STOaWe9ALmgCFr9tgHKyuWJ2UJ/yxdWcu4iMhZ4/8+d
QTxaxqjtXOWGp2QCT41KwyWyS07dpCZNoSA3PghpBfBLFtnVyicTg7UBZok/pq9P
vVgpIoQ4mcd7zMsTdtvstr1tUJveTJaaR6B/un/Miubpto+ZD+lpv4sBtZo54tGT
HodhOBot3CDb1Xzax7pu/4WL/jE7W47lM9mH6zMc+rC1NrldEXLlR7ekwp801fYg
mk0/IDYfwmi0vJA53E80sUqPvS7oX6PQw/MRJmRWF8h4lNYAm1l5e9w/+qYDtmE8
vwACKxnVJZyA6DDcVP9tdKOKUPUzdCNvRsDqo1c1FEgBf13r4+OFuIL3jGpIiEdK
d2UaaBntBZ+wQE7iUVw372R3NB0E9H8XtRoIDdjqc54elbBxYmk1ehr8BHCUwcm2
julhPsA3HSEiTM4H6emW7MxGPLWd9COuIXn36QQMNg38KUZ6ffXRbLQpeuGF3Ck3
Da8eh6tNjH9UWVLBAEnrk54yNNGSo0xabqAB0h95NpTeGFHXO1SoI2hjHgESWIJw
LuiTgrrdi2//SzBHLg1sT0AdkakSaEXIqkcqbJU4MAf7vJYWhIsPfJYeVA65GNqq
PlmLw4l1Wh0Ykk0DfQ4L7wFml6u9XaeNyaMKAGW+WmTIcsO9+NseOBJKGGhcaTes
ZJwAlhzEBq3VPLLJEjQUP9h4ysrDQFQ8IJ/J0d5wNQ0Ux12X7Y6TCapuU3rh8XXr
gV2IfZBeUudgntns6CmmjoxH9dykkjglKBKwBEwRwLojbYIYK0s5cPDBLcWpfVk1
1kV+OGc0oCTHWgtA2GLBsz5yES/TTvOZkk18V88UgHrUCQaiHGvWHUG4Qixdj47k
8DA3m9VqM4TG/6HqJMCvctQyAxTHbCQQ8gYiFQvslZlMFlaEu3S+pwzPfQ1l4EvP
OQmABpbG0AijrJGfFoIqWrDo6gYsJgYa8kqMelZUNrgyYd9DSvQD+Fghf7XEzsxd
Kbi14hD+PnjsY0XPCZf4hqGjD3R9A6k+7EhO6ZTSmX/5lLhEJEcma7OmHpvqlfHm
zLrHFYUDpg303z4pNrK1+eT/+P7G1v9xOOXmENURKta9pwlWj7i4NJIsbL6xQFUb
usvywtVLZPM8RYbNfeMOiE2tHMcK6HLU/iXxghasOFoiU3bYhmgKYxEBWAwjLhi3
gdLUWVcday7aqFzZwTOKojfkPblW9Vr7XSg2hFk3A5vKG+O1fh9EZWl9eIF+uoKp
dqH1M56M+VSA2CF8koRlonxWbAd7o/B9Yam9g2994RMrxqY444d3v4m6V4LictyZ
X1sMY9URF05dxBXOBqciZFSeKXOsTWhhlft/WyL7IdBgm466h+NhMUogB8iMhSvd
hIevpAwYFa1Piu4Xo8ahsmypqZObiX5LLNPxY1mxqOsunSFubSQro5L5ZzkwFUer
CU2keviZKSnS5eyzgl44cQc9hauMzJri45cLAnLC0JV2xFftoRWjaZMn72JZguZL
wRMdhSSPN+kV7OqM52/d2bYYEGxpqOxeky2Pgq3aSMkEF1WU8TRGeh43wuyBZkW9
tqRGH9gQlEB2WARGm0/osfYewYoJqLNJMfzWWXYD7wKZVjT3nicPlvE7OXlSKG6b
0v1XM0SrL2u9VqYcEc/MsM3ddtzacwzVzCLC9PQroj3p67lYyQXcmH7ue+Yaxsnz
7Eycyh+tKyCHsDqScYlpZDSHzpgh4CeX2LOUq5JIzOgcrhDSkLJWmgE9dGzCGg/U
HtqXrVqWEogGAofhHEMW1fZblV1FyHBPkdTxN+oDhqUYYkjICe3RKzDUQW5m5f3l
/FCm8xeRP+YgXvDsjqEpqcf/pSaxqdpJVV3VNo1vwLYJfqMLaV5ejum326vwOdhk
MwVzJHzVHLIoA9uLru71HOTiHuIogBkZcE3bQjTdnWviDz/GNY4y5XHwAYto22zA
akgDQaDjp/Ci1Z/ieSXvnvEGgHSFgxcHvxCShQroJo2jb4IuHKZysQ7YssR6m8DK
FLMgbWt+bSeBbWPOqg0PIzKoFqenbzUWuy532bRscTPU9vKXrWWnXNrRiWE756wj
wCJCdy+dlVZYf0p4eCNvXNf28D3FZWSI5uBSHY8MEGkbJGYmax7K7y2JiCHuiZSV
R5FpeOWZBmwtEBMlaxlwjGbJG7ZUaIe9fWcj6RjVLfZujhH6RpyX/iFRBXXv/PBO
LKhJenBNikU69wRo97gz0l9774l2po24YP0a8exC8AX7Uf1VIWBRS4vpS8MyO1ha
PsnmmmXbAEbFg1PNkKBJgZj79oihVuYauFOCuHgRf7AZJICJ6tXcT8Pljm6mfgCP
zi229nnb+ibnHCoC7H9BgU2DC1uRmiSoQdZN5qoFU+75jVUNnvYzm+FwYSOA4ATK
lhaPaswTCd6NyD48irCHED/DWul67zWSQluZi5vJiPWnagQL0TQP8GLqMDKkoTkQ
Bso+NAhbsYc1aUoBrXkO5GxCO56sL/rCCYNHZsQUpoWPyhZf9aZSJwoaAK2R81l7
VmaOuV7UNuGQB1uIb4o6XTUPsflQVGAgre53h/UTVazIYK0h8yh2eK3A3fz3tLO0
/oypfgaIgfOanRkr6NF1bzp4dXdIByUeeck97EvR1vgiP6xnJn5ePFkDeFh6SRvY
awWvL57F5qsyIqlFT3WTJJPBMyA8Z90exA6SKMQEP/sjbAnDemJk5RDvxGvf+fX7
27NQMTZ3S6EkqFaQJjkf+NW6Wgtt8fFrEH65diz1asH+blx0Lq2U3tk44RA1cv0G
wds593glO54j+iJpDG8oR/+Br3M+GsX1kNzdrT7fQzaEtCMR8AZRPKedhTftkuUi
XakHAbo2wt+gl7HhJUn+VeR973AftPIZs3D5M7dgeO3H8QUNvXY+obDpjReMZ+T1
f22qe37dSIeJkncBRfbuPnG3ofI7+Jv6Imsk7oSw+GXboa3InC1P7rQmHr9LkFD1
ExZDZWLstzaamqAgeclD8mC9RvU1CJljNAAHrtVHUDQyJe6UgMKc9C5+SJuIOOgL
uE6tCNmxdicjMWbRKtUkKR40w2ovgjETAgkuwEbmF9y8oyqYOcqFWFxASdQf1OHs
7CQ0Y/TLkU5w6tV9gLd49YE1kl+N1iJ0qTZgPX/OIqpYu3XdfYooEdH2qgUtGYRJ
HtDBAbtupKzOWaZXGirIBrxOIyUBT9iHyVFp0M3zIbNBMlFJLVRU1lCr6XCxOY/U
uocLlzUm61uPdolcxQbjMMJb5eFCHhmWEyM9RuQJrfsKjtKB16r5Sy3XUcyDIxUO
ZqATFO8nVo2sLhbDQq8O7t14F5aWdzv1SkFHhI6ZPKIzFMlXF3OKaRauQPddbFVC
RuGmNlZNfPM8zEUcHpGVblY9Q6Ntg6JyU5tw8bEx8zVDglV+pr0XOc6D5FMuzIZ1
emf0EujRIuFk3iy06qw8ZzAPFUTYquh+Cu+R5CmBcsgaS6OxwwHe2OaYtYZDYg05
iD6KBYkUeEuxoLLmQsz/dMyZY//tLLI3tWc41ThSYZohLAOExOALhJkz6Qg8eqTQ
1y0NHbFKidLghW08EtrxcPUhnJp0u81Dw7iaUwGDcpjjtLH7t3EXadtZH6UaDZJ5
3oEewkUoCi4lY7FWRL8crpBMJopeqfEz8FAR0a+XreJjcFABdU9G7xohp1JIZy/v
oiO0TY6XBSVwYLC/SRw0mgFI5trVIYDiGHhS8Adf8b+NHcbnKmzfQ/+9huKa3PCD
aKKk2rsvAOkDzD6SQUxb/Nm6rMeh21az2esgNZz0jhiJoY2S6LPWvrwnRznoi1Xh
npcJ56ccPAf/XDxsQ1cRR9AbpeVxiBkYuTA/jwFY/NQEOdvlwkYJuMIjPapENCi6
fk54TFAZfOI1r+oiI7OP4x9hS/cKE3euVg/+wyeJV75mHbUBNgUaUxLAuEeQTbJw
betXwACNbEzg+OK+HCy5O31tA6Gb6hvWGY3h5DCks1CSfa9ZYP9ihXdmXn4rLtZ4
KoRCdz0v12Znxu3i/KmH+TO44pjcFHJW93mbRkKkYjdpBf3yE+AzsBVUWASE9cqG
YaQx2i+TyRkjlptrIlfq2Kn5D6a3fKshspcj1beystU4AoWzDKo1FoqUGW9Yhxv4
Rpzeuoy/XA6fiV1PMHlUu4i/oAZEqWk16yLqoT4EnqIPQQJNk3eXLN82zOdeXd0z
VojIHpT2R30ilxGz7wFA5jA13Vf+aU107YpA5to9f05a5pF8e3bDG0hO4tMHZxaW
caMbbGKcljBCqdYIZ0Y6wlYGMUynv3wTvd6uOamLf0gFqgk95b5/DmzRBtNaryYx
/+PtKDXXkPs42s84qVrGXwc3KxiXSEqo6s8PeVBski82vFHPoDT8ONr7vMAyWIhV
6fmvKB63uVImra8AGURdInK7QtwTSGXV5vcb43KO1MWhAsKZUpmP5BWZjw1ckHJ2
WX+djPBbSvHxts7Xohuukr8JfD5O2ce91UBuOYOhsuElkdksaYLrxG0ovOmoliSO
I/8jtu/WZK3ulz9Rd8EchjM91m9SceY8uBgHJyIq4wNZS0zlH9xXLB5ineIUFo0g
IcBsgcRGJ1UndXsCCCDn+5qev8sboZQAFA1ekGvXYTea4X/QY/JfXbNxWJb095E2
qMNSjDkzVd5/0caoELFWVrDliboFQbX4gryIzooEVYuzRPRbZnmrWyH4TpWIBovM
yy482UmPmkOyyc5ZYklCJN9FK73iE5yvDJbFwwvDvya6oUtcwyxKszEjCc9v0aCH
1ZtCX3BJJIDWh7FRBEC8YuoUWMJaR2lZz0Ip+c5+St9XE3vmeDRS1J10RRL7kn5h
71Ois1AcOH6mZHi1zo7mV4xfOS6brGEOrpaFYlAe051dbL5mIr5rcMSz4mwa/bhI
0F8nuw09E7LhfLGHmDPpI9K7wgcNOGIlNwHZx+TIx3mTMfRLsMa2sjbZBcaS4GUg
f+txguPcRZHQ7iWQ5hwslGTGAIZt5ya/NRZpIZwSaYcRe4SStb+hlLOwuAOaVaQL
AEksO6tRuSgFkupdtoBmBPRqU8i42LfRzN5Fer+b3yf0b6xvEREGS2P74XRuuLJ3
PPHko07SulrG6KeOG+w6Uz4TW1bCily0F0bM8fJEyFNj88exdDW04BxIr6t4yFkK
7x6c1fWZREfgkBi9PXGNeiQcV25Y2YTkyMD8K3TIHNqQJbDecWVCtxy0mOVO5W4a
utXTu8G7HtJXL5uFJnjI0r9HF6K77aFQ73lyhWFEar9igc+GWA7AQ8hO0gG8AtMn
cQ8sMq2M+rheOqVyvcdrhhHAgo9bUo/fSaKWCz65CKWDzv84VcZcL9dqF3MjIQR0
Lk0xz9wlTqWJNPVNpG7yPVj4WzJ57KWtFrEXLQqtPIZMQl5vprXxzZ9Brjl+tSkE
mKiJAK2hVYTLDQ8s3fqw/wcCe5gG+5yrSiEvzcf6X5nohwonDCJelnYWBZ3midyP
WElV93j0skNW+XZVJZaiwUP36fziwI0yRLz4PEMtbTzoV6J7yTc9/cvYZtggph1y
AHfA6aZGTB0MfKJ4AW94tfxY2BdSF2b7r0Ok+ELhuLJk3RIcQDQ4k/98pHE4lHIp
l0w4AIh/eWBiROJcKwOP7vZt910AvwWxZSTtfAFdWdVnhKI/ekLxZK03uVCzopas
vgWbgvcdbqujbZAuR70AazgPBJDS3elrNQgMzQX2hmtoojUSs3gkZ+Uc2ZdUZEyI
YCbb4pq4P6TUl3aG/K8eZLJvcUccF0HEPomxIBLXyak6Hy26VjC/2nHzTDFCf5tY
/dTXvO2x7HFMrbUoMtbw/JmVfOfbmAWCW9yHg5Fv+GWnm/ees02ap28/GAoQ0kQq
sqoXi8HrkJRLZPg1OCp0wSkqyOx2vQPeXE7Qeb2yRLyrri5SXkOHFztzKqrx2DSP
b0G5lsZPw8zgq9w7bUvLiyIWjQtZIDZaVXC5eql+tmSboxwypWyFAYFK2E6izH8z
MR1Tn7BJjOsy3ozCM87VQF5df6WWdOkWlHB5HnkhItXwQSeqzWhbhoTCHQB7I6yq
p+3WXCct8+r2/FAl5ahyQa8s0FKAx+97gnvX8LundGCb4fuWXAEBhMwZhd0L/HJz
mVX4ZCafY5t3eaCH619MGMaqkmmrSKZ0duCgeeyx0V1NEGW6sC/GiqNfoXFzEAJi
8b8/ImwVYhfT4V06HBewYe7Z7IVM6VDvRw/MreQJmjhctzSkePgPh/8YvAf03m0S
lygwL+a852qw1iVzwaN9h3NDpf4KH7Pyeyr4aGs+3n4SZlfBaHTvu0cQoXx32wnj
YMWyydZRBgR1qYSB5pnO9g11x81lcVCl1dhhPVFaU4BwPq5m+LpJRRukxl7UXdJk
CSe/uChfv9y5ThhDIngtrx9OejW+tWGYCMnitYLQq+8rWC9Zn2WiNn2JFK/QYFy0
b9mFXO3O1KlNHGRf3yon7PcsxryuMybUOp8k4HbtUx54n1JcqPtYMnZcySQEuPUF
xQbYTaEAyaL9xgsEztTPlznou+XPR4fW8+p4qxOakRSMAr2lb3m55U82EJkj9fRt
HuiWdkIRYZ4nQKGI+5VN/b30CMnXqYyvxM/81SNbJmHVvkX6qKqHso1IoKzvhF25
uukVUWWdCvwYG7sBWgknzfT2B+TPIxfznKrVXrWtKRqrpiPPJhkPsa85n1FF/q96
kWx5515KiWSXaHKVDhK+cH8pnaUuqC7T7L/M2fxjQqvW123KF9aV4fVw4h4Mh+R8
f5QCK1hJlDhBxPE/mllpGJ+su/GCQ/GXvNyRYlRFO7ha0OoPhwUMenV0B/7kU2Kh
whqD+sMhJYaqhiBeUwjzyeM/77rqighfGA+COUId47MjlsJ5Qk3GiKui4Dl+H5gA
Bcbay/eSTocCxtVhKka3YcFVsR8egAnyHSSNm4kvytL4CiWfW+VRyDgMQMIzOFuO
SRilfFjoKrrI/oF0xDnQnTP6Tocfex/dWgHw73a9kcAK+eilaKodIVcEHsChho0Q
6NQJZndZ9g4beeFYjLi+o8bhq20QewogauBdLhaXP/g0d2OFSNf0hfj7kbNVrNbn
jhJdguS+Tj5lZgRs3h5kBWTMKycS/CdC8K7E69o5wyUFuaZHSq8a68lfP6T/1fHn
ANwbe25Pg9Nbv5aPk9ICQ0Der4SOhhF5PblDp/3gY2jaLkE/Ymx7W+h1dLQr7PPL
oPyyIi6MZZZNCkbXcY61OjqVFcYa74TCVw6gS650YFW+zLQrSJGaL8At/MClRgpr
hravFP+3ItbJf4tSFsGaRrnH5PMvTKMwrVwHsx/5eI1py8vS9I1hRNyA0vzDRzs/
886U0557TXbIQzinFTJ7hmJiXZu+r+O3ivlgls6p2hShro5mJjXLjtwpdK5F9R0G
maQnk/5+2zHEy5wgVe0lOnzBVRxT4IbdL8ACYpfi/m/gSyPj9XIEktpRTWiAg+nh
YxFmHxIE43JwipKvR+8i7tFxW1ODt5xP3m2thJOHBOnRcAfwRNvv72MRLQuXJZJ2
vST0BETEEVMCC3OhXao6p6YKfkO1kSCaR2Go4ibXtGmOwi8iLb6Jmok/rmqHYUhJ
vVoDZnGBL/1ZmTJl3IXF3tzVTj3FDpZXhPJAIdsXku3cHnZ0QRJ8DE3qPRGTpcr0
3u06ynJaB4PcgIJyCYQk2p1eYcnrNlluX2oFatz+ThSjbxWFn/CYgZbcMaHLGBVf
qf+5V1N0r6J6UUkpxEidxaoLwuUNoqhfZV1MvHNuSku/bc5NHCjVr/qvur9ohpfl
MPk0QatLIipaVNpvvGiih5qf5CSBT9TRuaCWgCql4DcvAz6hkiqyEbGFAan7iATo
BaaN2I5Rgswx/V8SmgYckCh1Q/YjGuyQy+Ds9vqTVK3kPt0ocgGwsAOs6Y7XGJ3T
5MKs7ZEOCa3ZzCyssLGFT6qNW+6165s/4yPicwH/NSvjVgvt4Dj6o3iazlbZck5R
WY3Zuw7msRVe1xvtPJjCpObS2ZginUElwblYNNh12kCXZuF7fsMVxT0S52PSmLfx
6OM+1qoMZlo5osHViqFkcJx69BWKoc78Q3HXfROjWmibfanHt2Rxk02HH8H4PmK1
kTG04X0JdkmckouuaCSiwoZ4MqGJe4+rhLiLsO6rj64HNPv2aVkgnRQ77P+ADoS8
KfXKmYI3EegCcXchx3QXJ/FdCC825iCEimLYu+lkNJ/iWuMaKaUgOGAEXDfdLeWo
lp7LWH7mTERJuR/9pjq5lnuk7hp7coLwAZ4WtZG9k7WaskCfuwejtBH0PwokemR1
Btjx8c2++Xv97w49U6b4PNZDLaNWET4YNrLclKaUTwTP8gBivG++odAUgUuc7n0n
7+qH33top/59qHP91pdsUQ3X/F2zc4ceLprZAtN6wea86DlTxYa7efB11Wh/rchD
KY3BOsM5ZLsMPuDjhECYhUKbu1seNexzUuWRdOCKzChv8I4SFEcbAF+1LOwsGsye
59CaOdraKJd4xN3F00+2q2E6g6CnQ528yWv08cPtF2DPIreIrIlQHrod6cLWV0sE
Azmtv03wNMggoIR54zNv+COLxGbf9LSSVy50b6JjtzSFe8ce1YXptTFd05Plbc7T
KBM1gLxY9H8YABd8yWVeaLOLNGYxobHO/dxx4QQFgo0/XrHCvew0CkJYWsyyc0Lz
p8W+XyP+rw1zyy7bsrq5Wch0Axw8XPSQGH/z0hI8M/1MBe2YR7ocaIDU9Snx+iyG
tC8kAukAimpCbqZeYhBZ/cKpe33Q7rW14F/9X5NqiKj5bcWkhoRChZqUs2Ks+Eev
ian4+M7SPkEx2giIzDxu6ElQ9ga6/UaTXpPcWBicDDrQP37o8ANxF2u1+Lpl7gPc
3XCa5qoJI+t4XBS9JalvJUobDqzChhQG5KfI1I1ZuN3ezjusUVH9aJkvrHrNcii8
oRlXgAWN3IvwNu8H1S64JzEcvlu9QPYDcP0ZMg+XBJggqaxvSvr6+q9fpiDBBFe9
ep5Xg8+PUpKdniLWCBr0x6nhmAA3TqRaqyU/YVxD225fKeVubbRk7uwTa4RzrwpU
x+R0YRFE5FoEGFmC5uPqO5zCIJpcIjUocWHoG7zhhu4u9gd/Zxb9jPmU6C79yo3I
H76P7gPJAn+MBbvbJoPKw1q46DTSEYHBIRxYOvO56tthnXyqexTEd/KjNcOUOZcu
awXLJQNKypYaHPAXYo58BOgSK6MfC2RR63dBn6pFjUnVaoUzCATgVrerUKIJ66NI
ACYvUCexMpL+WjqhM2JJYp7wyzWqJuG2rkbwqa8av1fIGseFAlFk2fZyiXlSKs+Z
PboOR3FiVssjIok5jgyDTXAiso5ull+HXFaoLKPPp0C1L8s8AubVqaTxUDePYGL2
SFmE6zNtPHa3JZk7qMTICWNi6yeJnyDHFmA+t/Yxg/HldmfqbTnIxPzMQ1KE8yyn
6pnHDeWIRJ+a/6ylfPYZ9S8W1kCiw11KyuLYO5V5OG6ZDmoL+e+wKW/7od6nosE5
irmT0CuGdvvb6r0UVh4M7yzJzPqiuBWcBcjmPTUhACHmr1S+qZPi/JKUjgjpgnMm
8Fv3C2ztOP9fx6KQ2+6N5Y8brXMZgqg6iDYO/4t/mNXpr874SfOCdtND1pGXrnR0
elqT96YhfzqvwMxAV7PBUNfccdHAK1QDiqXjSSibyOojFcrw08Bd7jwGMDoIVZ1m
pBTsZOcGLTkKteH2rQjRM2Flw1DEU+IaELgAnZI24iebJoH94OrN2kL7k0zko1i0
6DIggZxpizejZnQ4tqEsf0BsdKq1/2STxhBMFQfqqDWfbEx/3jIS976Ttqbk36WW
9oypZpnQE7SmE70TkXMyvBVXA+Ob+kXQ4xHrhLhDcD7QrxBDDEL5WhkeOemDxE1X
hqW9gs469rNTeMbsJHfn43yql/1dvLTfpZfBDdlGfYq+0GtZyJkRFV4ERiDX09zV
AYjlaxsIiieQWSLOj0yqSJyWmCYOaJfMQFxa8T2Dw2yd6AYbUE2s0fkZGafHhonn
Czll2pJeWnrk9mw+1zlLaL1kACtJtAvl5JESzEi3qgpmjS19DkwxRQMe6eBx9EC+
YXLdfE5BuWuTL5lKrSalTHPUdhgN/G83AkNhsrwTM46pZmPmxYFy9Vqx8CBiO1+T
s6IpYuCx0gjLYFW+k8SaNLbbF6iK2p2IYFm4DkRv6jR3Uws6Xjo177bdkQxJmDbG
LrQXKG+bamLRMcA/HMCt21MkkFxANH/vWLjjBSiaWCnYbknoWCbqnn7tz5Bwvip3
e0MtrlPVyrEj/wJ3iF5d3VnINMU1y+Hpa3RDOaf4fETI5nivVu/nfcR0gy5i2Hc0
hdVzuWoO/NcczN//2W/ae2OTigOKG4+O9zUW4eXpFSK+4qNDa4/yk4Vb6FwuIBsx
BU6nHvAaeAO93/3nyw70YvHqeSKf2YvqkvdAO6AHbX7SMaRPgIrUETrI4uOg08rO
L0tKmPfL6sWoNMaK73M+MZKDl+l/a+2qkd6S+QqB8Nn3pOor5iEDKQFqg8lGnUBG
1+slIq8qv6WKLrLx+HqAiH2xRwj46zygIWeGsTonDt7RNodU1g6aSs1mtsMAJFy3
ZRJZDqHb60MvBgtYeg07jzsHMYiD3f9xoWysHiBkxER0MaM7/NsC97hH90bnKjOh
J8VlpgmsoG/5MLC3ZSK9CNoMKNRSEIWVOHgt45iWAyP+GsuFn0fhXJe76lDbOVD6
MOZJxlsbR65kIy8ezMnLkzlVZEm/4UwBYKkeNto7V2+7ZwGDbQtEel3j3hRUEeoz
G1f5NXPZlVpGVO+wD/o7QoIIR97z26YxdrdP9RQGawtEeuvXeBJgdoV2hjDvsF7q
4RWMP/nb5Twm0u0CslGxywwv09s2tc2KB430lVuDdBKzP3SXk1V3QEEZDORlnrgx
VPO6Ivl35HE/o1y1oJzjK9jegAK2JupCifbf8eXpKkcthetZKfQl4rwcH6xyEYkD
Yq/6NkvugpZQu3iGsvWrB9l9deHn6b9Kaaz7Ewv6nBHQOTwwZ4B3uFPBbjmXmtNN
AW9jmD6bMe6uwPQS1tO1+yxOJ5/pFMLwv1x7X7prXmDx40xSv8rCr7wEOYNuvR9+
Rs49fJGaQQ0rxjDRI6cyYFm6qxZL/lCmQr2afa8hUiCNhc2lJl6AVqpeB62vBbtv
wgJmVfX9RkFTQVN0/ZD63UEOa13CcPmugm9UG70OqKuCDKn1oxWtskXOr0dOsT6d
8Zq3XZTnDSGgbsXVnI8mk+nP0fG9BCjtXBKwStHKBLNu+vxJ9+y8MZWU4WoZJbnM
hXcbTrKUz7gXCweoJlOwLB/4SnSxC6leMtAi12forPQ0EHHe3y0+83ZBY7Em5Lvm
PrsfEQSB3amQsH9Dpe1BEYJWhPUPQg5GSb0z02VXEYnWtT/IBYXnQMVnhwwl+TO/
qDGanpH8stxJUrRwcx4DXw7iOe4zGGl7k14N687Mw2xhVW3vgK/Rgc6G1zMI5+KQ
c1fYdZLbCXCCfUyuLcuwqZ0naadM9wWfnEKC9dB5iuW9B/q7kJ+qr9VqeSCdEQAh
qVzOBlxs0hF2NbA4YKyyFTWrcAqGTDWXLIhqH6sMKkGYQIDlTX1cLx3jMWvIbefU
SvGyBJmzve/nJQ1alFGXaOIIvBIRLGHh8NTspKqdZYTv1EnvZOBPWgYzF8UfeU6b
FOrSxInMc+mwHBPCXWcz8PzIYIb10vBpq5THFxnuejjCHKMI7TC4AXkHByKwL95U
aTYkT9ihNwxiThQMo6/TM41OyPEI62XLnKnvKqRTH4RDBdN9tIL2j6n0riT5OwcI
QWacOnMOCmt+7rrr5xTnUH+ZLqjzFvBsUGy4FvyRNX2AOv1o+9D3FwRejbNclfTV
gbbYeEUnN8YAPdbu4U4nPVGG5HU8V1dscYKLnBofRwJ21vAwnpqZHCz+cUE8JRg6
+5WItRarWQZDF1NlO95/Nu6DQNUOsh6LaLb1dd0Iln/Dj/OjL1NHeR2BUt218Gym
2cF1zKGJmruuZd8x6004q5+93mUMjlQMguj0rMJiUGiIOOOwRHFBjz1f/t/BE9Ig
xN8qBqFNTG9rzeRrw8uOEcTcLKCVxfMeez2NDuIc/h0YMrG7QqLHdZWXRW3Mpp5N
5c1bzmmiKey17U2T2LCxcRVLCC6+UMDo/X7U/VaLOK3all6pXmNgXL4Gq3prb9Hq
1B6FkNXDLDrZeIevbVqljBOO2bkP7PBTeWUNtyCwT+f3kG5wOXOCIMzG+tImzuhS
lMpUT8CduaBVwcSg5Ivcf4nztDhfXgtnz4zYHduaYxCYiKqosytI6+9CRwtFCxvz
emyqrAiFP81YQXXp1qCjCrsxyibZxTFC1s8F3JiqTFT1juzruA4cUuTE+0HnP5My
i/zlkQN997hJrq2sgP/rCwFaJXE0R9La85glgAWcBYjLTngVrNtydBqfWkdcOcvC
81k6SFvhYEe0VLh5fBMlxmqq6JkGWTw1rVN2MMP0cONwsuOMyYvXSHPNPvRy2U5z
dqe0aJstBgeK3gc4Kx3fNbncEFOy/WfwBt/1dJhLnsk4Pohy8tgydIF+izdfUgFR
8n7uN/tE80cSdePvkE9MB356D1skBRppKO+yTkS0SrdbIDKsPLKKQGduHUloV4Rn
8Ux842fnY8ZBLnoic2TyLSyuBk/UEp07+fcRR1KN8v9lhtBM635eTLvNTIjJZPLu
AXVKQM314Uslkv3PAdFtNEvxLmqbo2ypSroqg2fFunGsHwpttaZbH02k8wdjS3tl
J2hSP32oH4GXzPzIwp8lRirHNU3fQniOY7qFjAD3mzm/Rkm28NZvpZ62bOyVpS94
t7/lYWZWlW+qeo1WnQ2r6uUmrEbq2qdpTXdfLwUqGbjUstZRMg9oa5O+xXzpDH65
p4ZvShd68RZKxppuylj8Xxv+zqzR31u/mSklP9fN4sr/d7zNl8CcUaa8SNOd2D4W
KennURGiT3+nHx7tPCAp/hOFnCmwdmCaW2b0rkznyiQPLNXHbq2zVTJ8QOX6t4Sm
qT7/ZCnNkYaSKMWIlzC3cll1tKvB2aKYjEOh5/WW3K4HaRZstOvVY4ki9QWaVgcn
xHz61kUL7u3MUTCshLZzvLrsgx4vDZ1guWZqdXKSSWJBmcjNCOiU82z5OwGMGzC7
4I3IT8UbYVCrQjsqSQwEjUsxaLug7eoShGM1w/H/ydOz4m8DUFYHIfi/4mfsREm1
MjVYBf39uWN/0xdSoHvbtz3b+r6he7gO0cRSfW8ehIbmrprm2Vl/XRJLXWO4VT3P
Sq6UTcQMcgBgxyXX9VL67eicRZJYm+9uwUZMvGeo72TqvPyFmsxCO/NdIae5d91n
PF4IJl/frYiq8dmI6LM5B157E2CfEbBJ7x1NZ04FA5EF2K/w0S4xlUFWb7iwnSwi
l8r478TE6jjHi8z2acUPfXWk8yuZxEZNmO6XMbckHUJG6aYvvrzyoy2mG+O+2isP
EJ7qBPH8/V2NEGV6mM6czDzPYVZQfTcRcA/qMSVNvgSeqFoQy3/rQIUfAT0y8KJ4
cbCH6slXSBpRSFSWln8o3Xq198pM8B1Ax7ZAU3Y/8JAbcYxH6LpI2jwJBqPY8FAL
pfc6aEPaPdmNkivGTl6MFVdybMsgkNoteCVUYoWE/3DTTcZvHN5P338kIIVADHU3
fkFXICmv/rw7oLVsRqw+QsrphZ/uogIBhvTrJC03ux6vfcnZ7Cbhqbf16qBFBXMz
c3/nA7XRkaoR1DFgB8baywXGbWDy++W9X3hm6T/JgZCbZn3V3d2C3z3Wt66vNF0f
4SdpeIJAwCokcl26Q4HT5sRWyZ7ShYzbbq4m4YDOBaMetSuiq2Cv9a0ZMxRY4GVM
jKe0Aua4OSVjdDsMccQshv/CvOSIb2BH2W66JeX/FKjEx+1EB7Sfy/bSxc0HA5RY
02/dgJco+5FixXo3MPiiXnC81gy0ypeDgAoGDPkAwXPQiqom9qT1pH+OqVxC80SE
txkuKlpfGzWcyY2l6vgALgHyVyrZLOfXUjzVrGS3oVtHsJ4hM4T4Kwr5nr0ME1Zk
pIKEduIehkVG0/0krinaPVgycHaBJYyboj0sMoT2hzwib1bvQjvXu5D9UtuLIH1D
IemnIY8aP3fUvK7RMhRXQbRDrkmpFCKIV1lpyKYwixNk2v2hofkVHHcRZLVbw8Bh
/54ZjL4mGKc40k9qzyUcOAk5JIJiV9dAPUZStYBAIDr0rnnbOw/P7wj66Bslntx6
M8ewu19JVLarDK9CVeYnaIFRbkvQ5NuXDPkF43hnsEclbGRJyK+VBbXjrSDYvZLp
kOnptV5iebQtvPaKyBAJ9BUEakgSpX8lW9+8ASTnFD9AbtdWlXwwbwOXhXCXh2/x
R8IQ8fLSwXzwP6s+iqLUuRQij66waKh++QLrPLfpTkxO2KG9zJd48OHFZrTVmmI7
Pj+gsBFmzuFEgJDcpzQQvbvRdvOWT6+n63tBN77KKengDHD2PNoKbldDAeSuWst5
aPzOhdS51hX7RRPSgWF+GaPxVj8BS2hS+5A0gztGl+Zj4oY12OAz6G4J8aF+Mnrr
l0xMGR3GHqg5fJQcQyY6r6a6bpYM8AMoNUyGNlUiWjTTCq7qC3Jn9QZ4px+ZoHC1
SeWsgllINK9gFb4or7/alV2egYewWQ8YQFUoZEQPFdiPTSMhpuosfvkN0znly2Ft
77eI8Y8D2EEDa0lFh1GIB0scTDOfLbNRlBGo/erHpmLV1SivEOagHX6ZJ5m+rQRI
XP1RAVdFJv0kJVvf6xz3RsYT/l1ZNXTVoRnMl97ZvRS63Q6PaSZmt9Uf3vomYykT
CvecrFKX+23AShGj8Mtfo7kUSUUHFnGF9aqG5I+IBQbGsBR31OBojm8j6SYFekWk
wchylCdhsQaupQqBc18+o58FWtIP5Y0aUW14H9IBO9NbWn8h6jTe43c7YVZrEwlM
RqZsCjUtakFg/8qPhx9c55MKoq5TClbRMRDl6iNoV4fZFNGK0RsLaoG/mTBPNy2d
X+eTLyeMfTGwwtaTQK1wUqMggm5Wk9BgLbgVheJKc/7ZxMD7RV8fNeTm0bUttBoi
fb/LHof6/Mq6PCmeTfNqxLdsiKqqVBrdHaS/uslGqLSeKeWp5hfK49oJrOQAPyBv
XdQ3xLSpgbV22b5MjLlQoLmBFQwViFBFV2M3rjrecBIx8RMmxqqFYfWHLxxFODgV
fxLuWEW+T62gqV09X/rwaG/iS+Xs4qIxi67OWW2GElERNK+hTB+IFoX00+BBe0yC
CKy0CnbvqrXyzwTS+ftrbp8vTU9Vgv5tfLV4nxLKNrf7jM9oJ8v1qivmfMcCY38r
dK1CVhHshel+P1lPBQaxiCWHO2nn22Cy3amI/G4w21UEAlncui6fDVIH4iewthd9
UFRzn57WG9VXl+NHQfxRc8D8XJqScnaWNwqqMkkzV1IhiGQe0anuUK32AIifNLZB
drO2J/HS2qip7njKWcf0gYrSa9emon1/TG4FHQpnco9ofm+ANAe/EcIpXV4l2LBA
soVHsNre5piJBe6H6lBio4zHCi1igTwImITF3pKmorjm53nemshR2ZAgEUyROIkG
jFSSRAe+Ozrhhyy6Su0+jYo9agN4Rnm6isf/G9W7W39rBm0oGWP1YGgVGZ1H3UI6
jyKK1S9ybSCUFXqXSVEVfoNDh3E1zD6b6d3cEs6tgkZFEgRCPuXRxvg3V6BQddcC
AqDmIPwtHvRj0Rj6B0BySG3+lN5Nk3RtOle8Dkx2iwxBKbyP1g+Vb0aubxqXtTkQ
55XjXEoy24dfEdM9/1RXcTZDUmjrhWZxf3MhqkSYLwXAtOWjcZ/O1yC327uOFz73
YyNr0/kMgdRS85ka5n5h0LiVQnDP0o2Cd8QUFyShb5VNAdsm3SoG00cDQCUQyhYo
utNyqhCRJIlYNlwKXSuEq/hh7nF6lNcaFi8xT92ww7NetSeyMsTQyajcnjaKnn6z
Ayd9zh6+9WUBdTQVFHzKZQethtyTUySBYQFj5CQAbl9z/q5nrFy6FxwIgOEvAaxA
RQUKY7WnQARHpIsp4a0csaSrEw2+qaHQGbke82N7P/z++oxSCEpZrk/j8v8EQMCS
P5wxAPjaFmxAeUw2yNGocV5n6hVSocbaX1nVj2rjLM/pA30b+ZX/52svzKrkPW0U
ZuE5w467gHhycj8dif1zi2Pm1VnSQBtLWsELKAjlDN4/mlEuaayvzVK7t1Fk+sHr
52XLMsJNl2aYEPEcAcmJuhsHSgx/afboig41UiG5J9cB6ws68zhditz0BFwM89uj
Exv+DWJu82XWLXsRFN49U0DFVo8X0aXpykHXRUVFnXNL0/rV8Oeko7mUh0BoOSXm
Og+1UOb1h59wTBvkN6SNKBR2cq5KwmLuvjj6v80Ij8v3R6Peil3AxMUEtFhh19Dc
0NwfiBnYOvjohrrdDuuB68h/VmxJ1tKoXVnblPK6TCVKosQaz3a6yBf2A3QMsenc
rOYaYYjUrZF0//5Cv0ExqIXjxlBQJ508NcfxENI5Lfs4rCgN1OD8RV5KaenGKBBa
9kNnuEHzEdMduJOKa2e9oRF1zMg954C6W4Do+rM7pJevakdvdtZACo5B96stqxFv
h2SgWvipL7jUYhq1KKKwmQPpqm2eBaZbIjzTs+qsAAjL7fs/INBJaqGUm5hdR8CF
R6ufYnnkvy+awXJkLbDLUxnFJj/Y1oGrjm6y6P1/7jxQurjDwwOuJNCe/nvCO1vh
vni10TWpJaWA87XOv4Wufs/l7Mw2GbAYROf2ECd9/4VmnaPqhmXdSQgaf/dARiQA
mYQc49CzE6mRvRHxSa6QwPJ7Zqzd/1g1tswimg3XCFGaPlVdfSm3Es4hBcRtd9e6
f27h7si2mIqSdSGHs1y4AGYcjHVgGV4MHHkW2NVYYqwm0TDUWrAlXRdjP3fKPOLU
pnen4BW7PZoKO2043HcM5NsJNJpJqxo8QapcQ8zFMgmi7tZa/wTPV7EzSIkBtsZt
UJiGEmGTG4At+YtTcrBZZe4edY8OQjvehnM00GukR7yTg1y+dvWgBhgEA1ozuXUl
a/x/ZWMVghh8PfwFHeUJF/shb7fUE6dtX0FJuxG0xI92Q1eGBrdonkfhtuvl/nSc
652SPMgiliYPXZu3ffgvCZycC8tUW8jjG3XEw4+H0xsKldrenJViOS5HuZg1TPhq
MGJD4h9m/h0WlAwzGiQcPUDCr+1EsWq5YwbUkuviecjb4j5gBjG+oElUKGXFB4HI
1r/bB+lM/bOLavkswZng6O4T9XfTBJhRFmKKropXMhZwsMh2JoYAD/5eaSNFxyiX
JL4hG30S+ZYXqM+nwWue+bbRQmTU3SDcvhV/2PsAlNAS7oxBJdCJEucVyFJ29jqS
HJkeXGtWlwiNasCVG6NKn/Dj9UwXJDpoHpKFlBO3pqU0V9dA92rKeIrHS5N+X6wJ
T1VQ5kU2zZr+nq509MG2FA2XCiQSsoEyNeYdfDjA6ZKVwm/cCOj19XYJeHCIoxY7
Z6EBvdScdJN84Z5L7kihxeElqISFQXLmkKqsaLopKA/ACXz7LOwZE5GsgLmT9inT
/GtxwKgs1DOMG3HS3M1irQuODOI7afA1btwnohDGnVko1IfHBoftYeqH4L7/ny2u
kiRVUJlyb8Zw/JXIHDTtxS0kbUv7AlOsXOTzXLJG/08aMotYtnSHtHNQk+HHTYtG
hNj/adANV9X/VPYbx8L5n3BGHqN9wfTcZ9O2j3pMs1HhRUPJ2K/wzc4Z7p4jkpNA
z24TwsMNw+qVTtO/lGTwUf/PwLAnjycwiJu1Ck9AJ6CP3pItY9AKByszjptFNDCo
1OkPdeeTRJg9YblSwO9fAe2wbh6Ye0+1B3z/GQVSNZO+tHeWv270mXrTOet9Xa24
mYKW83KJ7VHlMlG7B4WdLh6/z5VObLOxQUE+h6UqGuV3sQvQiY6irGXr4FbnFlxT
6BhpndedXw20r44Svib7ahGma4+ql3k5cF8hkKXHBElro6psz1UcRrR/ctYh73jh
OFyjaz39/JJd5zsGF28+9VigZfOVBcfm4ZKnyRfyNZrB5XjylI9/n+vuOgptNkhX
d7qAJRw9zGw+HSpRwUB+td0QabFOh8MT745e9nHkpwotUv7d3cZUu4NxPCyVFRUS
1l+QOnA3jNn4Vfr4Z8XsAdxgo/zsRJlPfwBZSZd+551tmurQ+idT6yrQS7xusHOx
S6eeFJpDetOz3pMvapb4GLSBcQOyxnS+hSAHUNkX3s8/rEPqh1xN/EhU4of9y6Qa
T4wQC6mS6o1g/LXkr05PyFwcr0CgYxuzkSRVkmFzTMWlF0MHgJs2qN1i23QiopIj
Sprl8uBXTUI3S5s8XNGExGzrxL57gEBfr9AkUivq89CyLqwRcjYyaNr3qwSJX3Ub
KGbPItK2snGjygcneYBsKlZN1Kyikhv/+gYhRFiVdXiVvzqBcz8PLcd3WZlITkNt
hLNIxKIkggsUyoDiUkSBt/AKvzJGWdtMYIORt3DLRDfYwQgSqBe422hW21aldeCy
Dcfj4TglpID+RUAVjP0FFfHJV9aprTT9kNm+2497BvovRuMy7eabxJ00eo/x+Cp5
ChofJFH1z0LaP/eVS67K7mi1nwU+9fc90dddroxvcLAJ5jIEO6U4Hgs9ZMMaPJuh
7TC8hjAla1WqM9EG0Z9jcc+EaWp5bgkwY3nMO6Ya6aEgOq4hmB30v7+Che8M2qlZ
aVKJaTTjoEmRqnQvp0Q/A8K2ncvtruFY06YphIPTvGdWNWFEw5mTiDFck1gCKJIh
rgKoBOBPKqi829qdIQ8G4N9xrAF+SYmDdURzjP6agZoO+rprwWnKfwjcTfb9Xahp
THGhootVV/J7Uesj/jfzxdBwb3y647+NNr3IAaJzVX9Hk0VyuLUvUm83gtZBUref
smB/o2Z3L0+ZI7iOyh/qRPCICXyh846E3nvuxU0+Mkz++1ANKEBEt56KdECbROzS
y8EfqWseeobB+g3cQJFil/SQBmPliGtwKAaDxs9FyBLS+K1RZYynneGvjLnWBr3+
vT1lDOw6c0LuEDkdpqpyMZIoFALVQQGT0MlGV3JvCK75qMz5WL6bW6k9VsiGcA38
7j6MmUygbxUcGHE++4cmcRmVol/AOAY20YS5K1Ld2naOnIc5uWFzryLcQIFc5sXV
xh+L857WQlmycejR3zfBeOWMietNpOj+NAQIMZEiZBbUbX9waAoDZd7HgLPXD7m6
hNcw8+hXAXBJrtPXZnloxNZ/XlOYn62ORDADpKkdchqgqXSd65ACRTCC8dy+eGIf
bccDPwQH03PazzVDaFMzP7MOa0zTZIU+EnyHmcMp6AOL427Ui9q1hOrqaFg9sXeo
TGi1Xzo1N2Mit5EEDN0rya/Z4ZHg14N2Qa4MCXIKKOJLOCB10aNit76zEtUj48Fe
VAknvzK3vvKg97/UUT8ibL76XjllrbuRQqUnuvmXBeVukK4+4/VSq8E3p098Yq4f
+qb7+54MKBB7TAMVpmtaVlOgO8WqSWIY7iwu6shYJudGOhV7Ik+tL/mjcQ0za1Ly
WnEzQz8X2TnZb6ib2qCv1JF9Y4BK4Aq6DXIRl2UjDfkcP8yEW+/n18dd5GvObNA7
TL8eT9Gxq1Avh+6rxlKxve/UKs9ughOS8qi1e6Q7Eol5uaGr3bkXzXPo47A3UG+C
jXwb7z/P9QoyICT6N7oH+Tb8NOD86YFbpwxNYTC1hUO34N68FVV2wyB9R66678Nr
2NJMitKUHevPhwHltYtHWz3W42cs56FF78TMHlJt0rQBDKXzAhkS9M48YTdWystF
LZncPI2b3TZkVOJNTxBp3xqqgYKnPhEBIiVk/2msq/RPDfrtC87PhlAeBsBAI7XP
Ma4h/L7I+VBk2kgUbwekB3FB8U0CGtf8QWUEdh816P/xu6DOXl0wVSBbONeYTT1o
qBCpwYxh80se3EYOlAXgv4eyLv2eAtUelu0779Z/b4BznSdDXUTlub8nUwtvdh19
/VsM1FMwa8hZAusCEeAw0mafjqBxdN2RYP/aKSaw1YlEWyONFdOaq7r3Sc6CT0I+
/et5IFipE45tXjiuLbsI6lJ3jh7DO7sduaTTKvw4wMEEXoZZNextqaS3x37jF0ug
2e14GvJ0kr+I2hEzrihx/mHP8ASGvNFgQfvYEWzIlm62kM1+T7CaAS9XdM7aTdEc
nXWty2rbN1DOBiyoIs01BkCBm5IE73Uc5uJdgI38bijLQV7YfNAIeWA6vzvIMkOp
qcowUjMqm1dRl7HezBgfjXcyvMRLqfnF8ltPwnQkIQpBLQmpBCxiP32Bu6bi5RLw
39RqfCfPdkKzf7l12Tmb8bp/XBk+PQcHOpYDRoskGN8quEyOZyWdx0Q5H01rzq1A
BP8mjxmAyhfOIrujwmEJMHbTvlF1OZy3MMp8Az0mpEc9VEaCk3ISf2yk/Czy2yhr
xmHTTtZY+g4s917CCR4hFHpGZ6gYUUM2OgrXrAH/00zCHfP2CNL2r9c+aykgR/iv
o/L2uQnHB/TY8LoOvtFFQsE4GaOE4oJtcz7ndzqNZdmGlZNhETf9w/x/6ubb0/6U
k79c58VyDQlo4J4sGLBBLLjQwvFtxCfTzRBeWDy9hjP97ZMKlf2l6qjeAbJFDElP
+4+x/9BZp4+tfOCw4OcWeDiRy20+o/7pgIDhGZ35pjJwlFsNAe2e/cQKiuC8pcid
AW3AGKNRGmnljG8f4E5NQA/9Gsiiyap2ENd/DmiFOW0n7l3RvbMNBippny6+e9jk
Ib8SgWJIPpcgW7ps7/VnQSPTjbmqPtteDK80NK+y/SOXY2hCU5J0Kb/qAJvjeLfr
ipY8eS98Dpx5df0DTQZoUr7GyEZTbIkcmjnSUZujqpzfuWEk3lls2ymoSx9k8tII
+sYsMCCRlY/Hr9ysoz64xGut+0XKhVbnZshKjE6kBcZ0ovTVy32jmXwgQlx/c61p
WHcZ7Z6muZNPhSkZgd7eNcGBLA8o++PVgoBnGfir+SMukC58nLcO6Txkrza497MG
UDjWTTXmasgNxpYUe1/BXEEVmYPdP7EQeMU+VRssqoSF0BvrG77tjhWfCdtflp9r
CNOpi+oh22ih2HF+m3ANma7fdncmDMfVMf82icaX22tb4UkKEkzcfEZJ8dDM9dvs
PxaWpxvmAi/8BI91VU8P8/WAYD8V4L3/HzCCeyVfNiNWvULFOWCiV+XRjCTVz+uQ
7j8I8/85qkTJiZlFlDaK8VSxRofKASuRRPF7AFYEEr7Wo1qVICiLXoe4Yj5lGwaV
17o+g1hP/bAT32Sj06iFQa5cQO6ED4Nq8xxeM5dofUCb5A38Znm/B3Mq4SoxLRhH
NY9T+Sw5j5nlG2GtQ+mVIREDsi62mexCtC8plfLqhanAB3ynzUl9A1n29/jQl+Tm
l89iFErVWGyiqi48UlUn3FGpZYffO1MmOT5xAEbbloYxzHulUW7tH+S1YJ68QCHs
YaF4s0/F3XL50/7rsWJsgCQmQa9bUjtUKGu5WxEeFrss5ik++uq3WbK2ZtUxWkgR
EPhfJ9Dy4pwQZXk7dnVH2T80BYCX/3+bL0nEDj0TYNFuDxhvyJey4XRhW+nEIoAV
HFHLUJSJnM8GHU1iqwdYKbre+kZD7MVeR8Oepn84pKu3cE4jM8tyGBmziPfTHDcr
8jjkrNTFHgshSt700uXvbH2pJp8U51mz3FTl/vMKuTz7M4lBMsft4aci8tKiJs24
WsnvSkMbOXEZZ7zcPJVUXkgLU9Ps5q6EzGBa03VSm3BKM0/RfzTMcl+tWYwUZTzd
4a25j6M4ZIJzEkMt1of8tboChenwZjxqfMDnIT3ltYIYM+IBgyPtpuUrZiUo+KB0
ajvQG3wmEM5Td4xpjYXARdFGXy7naavvgMW5oCoG0oh2RnLjKx7t/6vRxtuJthU9
lFIm1FKML1B7ozNILbJqsUx3LFZOGKwox3bWO2ojTn+KNH4jWG5yfLoB6GBDvF4f
ZJj838Ohv82gjAor4SYnQVk+FSTAjvw4TCz0Ky2Xqr6sgWiMZjaEQeicxoRHpOKR
TYQWTOYOejYiv2YZMXY/838yssu1k+QVnFbv9Pj9gB6BK7z15y6ZKFmmXsBLcab9
NBD8EEmtCvUQyKV1BQuloBZm7jNuK1N6mESVI7UEUKei2sDNd0+Jyl/rzrCuRBXI
xli4lzmdmXGGawHi+G8Awoyv63COmhnEoowa/sOCW/U35IbXGu2EgyGlOzclEOEd
LO97PU6ULG+uQiZKdaqlchgDIHOkVKjY8MgHfvMD+6BDHsZSTIj6pdFqw4FgvpLI
KlkTs3T3312ITDAZg2Ll/dWC45k/uGtph8oTPG0ByOpqgggN5F0Qw76QOqVnY4la
rQcd4SdAzXbGfTOcK8KM/a3xZOfn4IybEYQOqcPRdok2XKsMsSPMpt0g23mIGWrI
yV5h5bAHetIZy0rBiU4OGfPsC4pEV/NLF6bZXiDccrezde9qNed+BaG78d0jtOFX
/vp0md/C0cjfW4VoSGWiLomQiN/dHvSmRxrBfSgIhUIMy7SkJLSau8Jcoa6vqYP+
mSIwHoiTARbP3byZzgeKKA9xZeJ8+AVljJ/akBz8U2ET2D0NoDB4kXY9cNCYK76n
tV/TnMXTB9JNw1d/qOPvZl6rKMgoUeFBPSP6+NyGSMDYJpR23YC3Nv5mtRQRmfDm
p9b0CixElOzcxIQFIS72UH2i41knuqM8rwLLow8tmfl0VMV6DYl3UeTXVCsE28RZ
MIoJA6uRiTDsVL38/jOsmi3lFdRchoCpmOJbYaZgIk2MYeKkfN1o0zjMona7KQqf
qLT4bySszjy04L/wCbxm8y/BrWPZbKjat9VvTcAZpAHMPIciZO0OZfxU2lU4snOB
B6tUp9BEgvx0E1cp1uopoalWTAmu/T/kUWKmOuvNpsTWEKOAZIpC+jjn6MeKg9bl
fdmtLIwUQ7ZoG7GwV3pX5tdaxIgKJfQVs7mtP81K8oCxdfN5evGQ4eh1BsCLfro+
UaOjPKQSgGiQnqZiq58JU9Mr8rk4fnJK0aOby+gNKBUawTWScjGoZA+/aiOgaLX1
LI0XLFE/Aw61JUg4KqTPMzKbxsSsPlgFop1AKFWExtVwlVZgY/3SVW+gVA/teeDE
whWUwYjHhcMrHCgMcRqI/wIPUbuxK9ATYhPkgvp5xh6zsz98TEyWOnHof3D3urnj
il+WltNn7kolZB6+xL5vEhrZ2+bY3jdNqGBaeoPrW0rCL3B0lzA7M3VNBF2tcIyt
wASpI1r4TRdgyvSCCbwsbnAHJ8Bj0MssGBZJHnC/QuYcJ0TcbV69lgMVpdPARnyp
vEWfluu+SlK5peAfPLYDpntSgOatWzRdXXjnC+QR4Yfr2+hQsp1VnUH8uTlHeKXB
2ACYJmQL8aeqYMN30BqOjyl6M5ftrGR6gsgbxbeBBr6OR8yPR03ZwJIBkLe7iS1i
NmUXt+hopVdxyY/yO+B2Q0l28zYAa5r111vuK8GaVzNwd2bUdY1k/DBsS6HZ2ZV7
w5zhfLub/mr97G0Af0j7BZGuT89fj7tYclurn/z+AHWEZvn7EWh2V+eqGoRVnU+0
/mnGKBzNklnT/4EqJWp9reVjcVJBdVi5KrG52qW9HV8kNf8+mLo4Fsjt3VBXaR3z
WO99KOXr1yXwdZ9yqwAy1K7n++xqxqogZPJevU58B6UqdaCrx12Uz04ZzalNRILl
tHapMZ97qfNzIhm/2hVBDa6qsobYK4F05lkqpUwXn3l2iJsALwwJknLDc/YwcSf2
MnzDjbNJo5KkPtCOxjjQDgIpC5LMzz3YBl07ptVTt07rX/vunnWSbb/Nj9mI7xZX
j0dUcklanSGsN/BH4k71aqxyAztBsI4cB5Wu3///mLgCzM6kYVfnVYkFzPlVx9Hm
2sPiBZz5JXua6xZ1UZjCciL3YPuEyYfTp8BCHFlka/9U7uB+a7mZ5tV2WQuxS0VV
NOUdUrVEh/KrAEwmW9RcCR8Oyqk8pxO5MkVnGcL4rIpB6zGhCuXF76DlOh3TJ8Fd
e1PI5vfofwOe2mPRyOfFvl2zPAAN6+oS5AOyfJgZpIazvGJDt6vDv3c4wrRUepdv
U/7Sxtk2fEp78am/MjzUmddZHRqdhgfEUhjZiqMaWQeCZcyueBcDbn7CGci2OfBF
FswIHfeAKns28U5F5ro4qUGMaaqbYakxUHmI8HSYzvhcJHChA/AqJJZEaMNlSpTu
55I7YnJP53ymVHMbgTzTRFbzjD3PjeIGhmq5rZHxbFi80oQBUe2Vj89HoT/Vy35t
Ilrwo+K6ptqsctjSHQ2k0fGa/3ny1C0i+4Jg08UarIr/LFDypZwMYLV5QcnnTNTy
524jR0is21FIPHuyzD8EzwM/xCzYFipX/cGFfCEYqrCPC/+OyCJ94iTILdPnpqUU
A10dugfKReOHHtpQA+FicftpMKdBPetnicpbByKalclt3gRUkGfkvJNo1ur5Ksl3
kOKDp+nMr8P3xaDuvhA8m5OOj4nqgIAbqO1QiWghXHdq9+xDDYhypU9RbUo89qpB
i5Al8ANKVm8WyPvGBbUrdbdfGcVx5eaz4g/XMmACHkOApgM5arcBwGnOV9TV1ZUG
3i7cInW2NHUHxvOr2zMpO1kGbXojO43KLVnUwLHcHmoKESpwotSknWPzBHicBSxV
LgPK6mNWJrogihfoQVzv9ARLysZQq6AubLbkMjGpcLZlAAL/U+dBOk6YPSjUWysS
m8uBFlO88KG8AFUi5uBJ2TMYPUuT54mLTu6JTcxww8YhrfCQk6dAALBvQ5IRMIlx
N6NbtAfAQ2SjSz9m2e1RZ/7jBJxnbCOG5NpCJY48mmb3MKmRENTaBNdLWSIc6mOD
6TjjT72c10sB3JKRTdxbGumludYnaigERNKu5RSUI1jOT7Bmy0e4RUsP9uBYKyH6
W0SF4Q+8NHWB1I5qDqfvFGz77jCpWOsc4bI/UU/ZVt+V2SR4ghIG2fsG9rbq45C+
RftbiEk6NyIR5qr7bIgOeocdy6pPk2ClorcX18UMcIT5cRZa9jwQbdXQPES6Ah5O
v/8yD0CPoG0/Wsc7CQSl02weL1haL7suKREinWS0I0Fl1sGOkrL4j/e1anvP/+Nc
f8kC+uheE4ihCy3P4gLkCw1NkWJUed43l+C/UTVTuFMaueXiHmFebBFhC0GJqWHk
lOHkxJxuDlAQ0AvjSBuZse9FCbRr0pgwBt16YDZPN7GrXPZ6kXB4dKtwUWYdhFYo
hJD22T3N6Bd39iiXIhySf8B1+TiL0sIXMcabAtNehpCVH5XLkX0pp35ZJ41tbbaB
s8NK7jKKUL+m3RKz3+t1Gn2W+jdIJxenytw9joFMqbquxnrRDYVsBvdIx7wCjqQf
zBI8Uw1xyR5d0AeBmROEL+/dKw0vlMkfmNpcZ/so0RfexiCGtpcUwyGYOwjoUeH/
rnzO17dq5Oajgco6WhWU7Cb3iw7zU/jRurIx1+XwFhuhXhmtCEY2kSg4kGEqCwkx
VOTwhkGIdVbn+ezzGZF2AVxPJpqclNhQrnw1yogh88j9FC34vHu9CfqTjqbXyMGo
Efs+0cXPl9j36/51OYzLre1cEvfk/hcM/0W5mGy8hsFd6GTyy9WsiypJQ5JzY8Rb
I9oP/DIlCtVh1kob3EOsGEXUNpbL/0j6LiCeNmJnUFaxwOAc7XNBWi4Z7XBk1bfG
5QG8GVl5p0tWer3KRkna/QiX3Rh3iWfDKVhfFAdI+Yl5V4+wgzbD04LJS6SAQcsr
0ogtMMbpR1mVfHsAQnneZDBf+pkUYhUEfHPHUZS79sJjU4uqZCCcuf5NLN/WHgB6
nnw1bPFPrB/9FSukX4oUPV6CUVFH/4gXOyB4MeQt6JdZodOj2s1Jdv9mYN+08mEb
jEN8TWtxqMnLVqF7d2SLpVlmV7P3GKbmSGWXZ+bQWVOvLnwZvALRYFLZRHhx4Tt9
BVuqZSevdXwgmqLFySv5/2A8/3g4PsoLpZDZ9JLUjP/I9Vi7ZzU/UHMm77gXteOg
3dKBiX6z20fxm5brCcTkCh65a12dRon5AMHMgtZKyWi8sREiQMBDNSowUqNrdthJ
IPn7EgFJbBOL2144L/TvStHyRBYGz4wh6xcWaiodFrQbKJOZ2LF0ImZAvd2IaACy
Pvy7+C0ZdIddayyv71VRLr6HIKD9Ixa+s44XAJQ8bJTod/lAo+EfR/bIgY1J2TdO
6VEG0GEYyTJq7pgqpIjbcVToedcIsB1W9kXgBMIrkV3vaEwTwi/s8WDqioL8ozTQ
X9qoVomb9yMWuA1W4ZcXET3OTM94fcwWNaMrr18QqcjEKeBCXpxD+BOG0BM2Cw2m
i2DGa109zfLZvnzm8/chtakABDflZQjwg83njCrpH+BLqK9PPnHLgEUISxYJ/Vif
TTUUcwFU9BMh9zm3X3RWnFPhGJboIoAgtG1wZCA7g6Aoun8qwXnceao4nYeb0PAh
Ztn7ufi1gZpDtfOujBfodwBt2Tl94KQZiX+pRWYSrey2BKvHiCM+KZyL1Tao+/DA
zc9xgtWgyF7hdxPwxyd7NIY6r3nT11IHD9zVepetxTHSEr7OekUfC3Xit8KPwY0S
WItSe8rHDvmpT3rWR5X8fD0W54FeAwkK4Q6kVYTLwI0UvaCS5tcHDhjakq0yDJ9G
5uKR5IrT7bBlBN7axGulIBaOOAqtTDgoaUPaeZPhYrlh8PySh2NbQNGRIPaO5B9Y
2gi0v0jeV3QFvYzh1MW96wlDvGG9XSkQqtUqzCelcrBwKtxZXPNfK29a+ZJGJdzs
d+7YocLfEx5I7OIfoJblEIcxu/AoOT/wR34B3PVse/Z9BbjG+bYsonZ8CbJS8KXh
WCriaVSeCgAlo2+kHaCuo31sx/v0aF4SMo0UVnCH6cSP7xMR8sDvFFuZJ+FtmQJ9
4fNa4srT5Wmye6rBOIY2hcDeYZeNET++vmLErfWS8adB5b1INNLkl5hOcjkXFOGg
X3MN8cYDF5jXrwKBo5+nXEdDbaAhW6xQ5+4NWqEkTlJiTEDXgtr40ygwai8e0T8E
H2YhEfQX01VxhFYUX+og0VYv+S+/D3o4/eoOkC2BvVwBGdtgugd+gDAaKesBjb+t
MqNMqVR9ygp00mVec56R9f65g+vip9TE0wa8Ol8alks8rHpxOGRBH4FplklFxtQj
vwKodSdunqljC4+dsgP3tobX5VAPQwFBNlJTKZZk0N3JJq/g3yELeirx5aSGk0dl
00gXLB8xsJJ3ZGvrbMoDaOR6AMmc0+LwzDfirLXnfdF4h0SpjEyl/juItZM/vxe5
fduPlhtjqV0DFByXLHg+RJ2I5uf96VUT/d6Xwdrie6EHx/YVRo2a/b+l0lqGlo6u
WDGgdNfyWXH1MhEW/tFLYhCwGLQ/S6eboERwA2+87jd3wZRkDNGtVREfgV4ftbAe
6ICNsAVjgQZMNn8YwuEGQXP4v6jOoBCtWNgTfkBWM2MtzHIXSlwbcpdckqDiQL9j
QxAbOwOpVdT4qZZdhu0xcfzUT4dwaTV7e9Onx/WrJFNHfcpeOe7ABtlgepa8IOmq
ZdmX6J0lLCAeOgrNZBamEctzff9Mqif4oG/JU4xyijJho6NsILhdLnpa2SV/+dlY
VP9x7kSR/cqGkn2CUZug7UklX+OplrfJp4BtOAJO/vkdNGO+4xpJh6RIOsgSa8e7
9yAaB9aTiqcdb3IB17roFJhP/zWY4Qh85qhV/p3Y9NQGTCh2Mm2lSSZFUPUpd6c6
d7BY4GNNihNwvxBLkKYzE0sG4G4V/4nRwOy3Nxx5WAAZsrnFLY5t2OoqvKH40FbU
rrfW3Z6xiMIfPDL1LNIANt4jXvnNIjB6gqz9Dm/g4MFM6BCq8OGyJ/kpFtIEuuin
dC/8/3PIcn1WtQ5TsujcIJeOQm63ZpgoSDV0nX9nxa6WfXzDwBCoKgzeQc+B3jkl
tlKLzM7UeSIsi9WHRgaVj92JKbPy8/FPTBEJBnoa8AKOE361FssTcGBghghIiWWG
BHFpA/OSNLsbAE2ZxESiQIxy7SvHgBSUL9Oskn3VtRZiQ60WyFfO8Okz/z+fSbLt
XhZJWG3eRy23fez6jdXMOCt4PdgFuy250T2+guIwDMz/fksEu+kxmPO7OsZLWEnG
+E1TsW8xXUFNa3FqyenuJDRXat44IxzTSGofj1SLcKS8QatyJzpyFkH4VKU7cuJH
LN8T9/UXxVW+JHBmzQPUYaPWK27lNXwUg2HhZM2Uy3zf7XvNrXFq68lK2rRPhffN
Cjp9KlhfhAq3/NVW1GF1SXY+nUaKmPGHtacPr8BIV0HbhI665r1hGpxQcjONR6S6
GoP1rB10fyH7uIyOYxO66CTPf/I8RZfkM6qzUTiCB2/XKpx5L1yPlsxbn7rsOGHE
f8VtdrvhyMY3hqYgVaf8FeB8EQ2GN8SgEKPig/aH4kUOH1wonZwMV7dOkAU6ESrp
hnaMqN74g+W+h5IFgATAFSEC7IR8TlYYw6lkw75rRty1YRMN6hT/wBOGNURQ84j2
gx8qfU6j+t3vMUjqWQ/FG0p/0xBeojIuY4w7LD2J+wpHcuvmzii+nlPCcTLee5SY
bWukcYy+DOclFiiMXL30zQ379ATWm4KTuYyqcAIWtqUSSzlpJg250/fpUH5P4D6S
We1T4eICiSt9xtCzE1FmE47B7Kg3wOLkD2OhrBYDFW3F8RXh0Ge5Qfio3sj75788
HhEIWmXYP2rZmNHqHVgscRBSoShC7P1T12JBPAqJOms8RMy5bpWjnmipafTellds
HD4WoX8SWaYbm26hK0xFGjz498WKC3DojXVks4wx1j8SH4zzb0qzFH5996oY3/P3
buOZmChmmAPqwsv3ku8dBTxFGEZnIrGy27bu6A2nnUV1jcG9LO3EBqIWJkoHEpPu
+Gp8tql4GI1HUhxXixjmNZtKNI6MDl7L2EU/n+xG8NatK7zKzSVg7ou/6fcGlgYn
6XigqW6VVd84cM+Q0W+4CieBFiGVzNMlsGV8wTx803CLR7r5oTdwlOLlE6NjgUJk
2adT04IbubOuYhQOJVgM3L2avuGFuy+7WzvoyKA+KBvg5GyJKcCQFUgOFRxL6AAh
erUEklko0U8r2ExCDVSbNhKqjmD+Pi45pv94bZPiGwlPbKZU8BFlMkbB4jedPedA
nrgGNd7h39Xq0lL65SvFYGs0FG7i0Ke1E4Dhe91mQmQv211iWj7EFsp4uQGViPPq
kB7GS0FbtRZh46ADCEIOoSWPrvTvB9Nd4wIsPTUdI8crczMB15ESWWRHtcpITRsn
JC0OaGCXcHRtb6zrMTAhoc84Zd16DMhMh35C27eEAwMMI44EBDDqD6VBuixP/h/8
MqcW0t0WVC1y2Vr39XLeRy0bBU+VFGGUSyIiqfONAWLtOzvuPeeh3cHU7kUprDHo
OJj5owxkRllCal2Rj5+YK0ueYaQT0N+0ewzErsURncP5m93TXIxg8GLNbADYx6iJ
JFq2mzMaN9qv+dbbo679ozEiL8itdm8YTW17GU2YXMnzeNPfe+5GlAHbJxtHTVFC
JNAIH9fLtAvFExWDFlmCMvzNqN+rfE3eeexOadETDFPglGpI2l9ru8efegD4EYrM
B3fAjGvJ2HjY6oyw/KauuiWTvZfTEk9O3CszkxYHjAUWQrkYDqQ35jXsUQftciqy
XKF0DNY98yJEAW4lfDZaaGuCHxDkzlegzZjrBpLcpNcRLBfugLpcLlbkQeP30Voh
4G7R2vii/HI5YSRLmp5AHIR0TcYTFvbqVWWY0gC+kaD5K+gKDt21q+IvjV5p02cX
7uvg66Mu7+uKOV2o86299vmO+hJCH9efITnE0fjEKi0UwOdO9AZhhyuIqv4iGtj3
Ugrayz5DsCBczWyopRnwJVDynUTQ2WoWy3i8Fj3Htl1wux4RYistbTLqHjHEpi0u
Y+fd6n0tBY/Rufxk2ytQhdHFFWuP8tlc6lKSrJb8+pvl1o2Zm51AuNh6VSjd9Oz8
Za+dx8UXyTUdvH6/s8KqcHZM0D4uKqIhMmt2BvfGkXxttIsi1dYfpsULqLoLzMTY
XBpkxDj4lUHOIpwhM5lfem5C7zlq1BgG3xHqTcJWqAeR23q71Bd8iHPsDQlFmFlz
xcG6oYw/DgGKMs7zGOZiomGd/oLMKFugCW/+J3bKCm3S++WiFqvq+8kkxQhlqVr6
xZUTdD3JGVKtiUmTh6l0iDF0EcJN8EqPA6IuduLFA3mi0ttfhC69Im0+20cmGrYr
bG+OQ0zlLzAKmc22BTED6gKoZkUw4cjbZBViDCornAOgi8m/kp1gnAO6OFmbmOiw
ZniRJw3zO4goWIWlyUyieqA/BKcSGkddYc2zv9iRZrh+yiFCEq1uUyStPY68byMu
e8Xpe4ZTSxLgtNLY9H4RumzKCG5o/otiLCLIfg9SCxa7PZiv8wTM9DXtAkuG4oUu
RZWUG0S/l7w93dQAYFmDqSTrmsLCzTkFkJUSYGQGH3DykXYHXH5TXHt/e/w/Q/5e
SrEHHF5zLreVe/GNtp8B1L1A9kq0oQxMCmW9KHMFWf9p8KH/JtRvOXrF0dp1RDxE
21IICV1FFiERFPQILIGRKmsm3lIe5tpTccgf31OldhT+VB+C7ucVAdlu4p2BwuB7
pKlLK6lrZFNk3nE5IFiGitSjcmtGFQxit4+zUlzA4qh7mbnoKjrdAj/gey7KcwOI
mA383EPrA33n+ylvW08zGDx0Rz/ylq7hMKBV9u95gCPmDIohle0aw5s5t7NAGPlp
Lsqcca+cFRnBMLJvmTnz7GGFkqgtd4cGcINBKk8w5ZAXAhj8OyHPuzmCSJfBv54k
kpVj4vSxjZGaU2Y1LGfZz00XTOip5IyC28U0Q1H9t/niLIqmPGeFMTVwyUI9AuyE
Lo2sEwGdf4MkpnD6gDKpdL6U8ktbPk+bwxYDimoSmFARVThC0P//9A5Ir2jEU/E4
74kyVzrOBdPUSO8ts6d8tltNiqaW6r1NDw2l8xmnmduViA3vTCYYvpUCJj5zFs7q
5gRVczkcTvtIv5RRxbo55lBsg19ihetuTHJOyafyxx2kvP7zV7aZHBrwTplmaQ3f
Ce2KdTg/9NM4RhDJyP744M0XYdW43sl1zHTgxV3CbBcISdDiPVvBD70J7sXnJrb7
FC5ZzUOdHM6OuBqCYtnTJzkiz+zzZLv+Abg0aBNT2CW9d9PsdbiZkcIdlxrk24we
L1UFxIYyMkLvSCFV6wxOH+EcOFV0Jw6VEUEdCi8RGM7vz0aw0v2poXwhfs2nq2Qe
JK/QyNp/Z1CSptZyMuMfyjrrRmEsKHcVvHePzU9p4yhMkgxYcTUABWFmbgyk/ubr
5RQgBVVT++xYM2LcGG7C8fDRdS4PAHcmyVYlsQNatXWnzcHQ8UKk+SA0tWR9wc9h
QQROWUoIiPhIrsU5Op4v3mYvAE902hCL9LW6msCuEVNi31buP6HirlHMe/lSFiZ7
ipTEvZJPzI3WdP6ikpqxtzuJIpHgGfGBSXR/1Vi9uicwASpbcYsmMNbICvB1BoUg
P5Lk6I7o6WuOQTi4THw91jtlh+Flogtitym8QpqqTsRkKjCCbXMVFdownAT2cfGt
Fh3TJ0GqNUehFygEGfalaEae8S/OYVTiQS14OawGf0caMvCGcvXhBjsU7IywHGek
BsrYYFvx5rw4mWQvkUy0tnWy/lxh0dIlmDBmc4eHDRNgG+OBHox2Wb8S5vHiVKP5
DJB8iGEomUs5OUXEf52mof82kuz2AXW0BTenBlq0IUM1andqmIJkZvPBlKLknZRo
lZPn65ds7j6zsYcZlEsGsGOenQA6cOzk+jHe8m7AsubcVHX4f0ehhTomp8GXVUKG
IKGDzXkGlmJc6AkZ08QZCm/v8goIpfIu4Ro1L4C2Tg1XqQjWDwudPFviCpVB0R4v
oiGmQ/nCeokHn59Lt/d2MsJ5/xa6qs8D3OPVtMxDlT5IuWDUErTo8TEnsgG5zD81
CM/3x60OPp6uGQQ9SIltSrNid4xjNNtILx0/jMR2yMflxJTi+MIfozdFdGTEpIae
ePG6m+qZ0Xhqoqo7lP28oMfsbrW8Qfy5DICitM6dUj2r+kC/EzfGfO0qbZOxjqo+
HoBSru0qlRJRBQgmYR4GBbILyy4ABQQnZy00WG2T+5osXe3YLiH58DfNR+Un1x1j
Z46DD7SNEVuD79vXqSkVcnqEt1xUZSHEHIF6jzA7jeVoSNIIU0fJA6DDwOa1Vrzs
D6neWQAKhUi/sIsdwRdHky1mDXeaTGyz04a2vRXkBZ1DboV/hIj3aAf0nixg55iH
c5hgFuaoHx/rOFOfVm2u6EzjNY13sv7nav9v6mg8jaRO+tg7PaGeJ0r5YS0Z8/vY
dMTlXNDLddD2zFm0Dk73guB98KtjEimh3Ctd+lixZJUfSD7PfFvG3zzGnN7wDiOg
TfD0wtlr8uqVwgHByLihgqgsV+6Aj8oByHjRhSHQbCPZOzqvWpVdQFpynxz8tg6w
wCZRh0ALRTB7Phq+zrgOFUGATac1FH2BxKMYo/0shcjWOVRJhX6uPz/g0u4N7ARK
OVj0QUsJ8hmxX5QP7KFbG/ighLvW59OYv//cblSg9YJHT8YJmxSCBlq3s6QJoSR5
xVxlrFERS5Fjc8hDsVDWqqu399peoyBRMsrq++n6Xh0jA5VIb6ry8CcwLjZYGTwu
tslP9yICBGLr94PGqoZkZFFWyk5NvaZ0nmT31u+w8AmgZBh74PVLbaj/iH9kUjnz
NG1GKLDq+9KJ1/cqoIbEknlcFlbxbWbxYkRBGfYtrNFwBSYlC8O+Wt2Kg94Bqh4m
YobHctg/CgQZx7TV3oKJJNbbT+XiozlPJjQyXQxvhnh1buXz9ppjIcIIWrB2feTz
6AYrSadnaw9/sNwM1XcL4OvCstgsJWcqGgf3bwF9LDTzdR3NtVDEiUjMJZmTgY6V
EW3qydkyRbyUyMFULA31rRIgyQZnEPp3z3f6w5YZ3R26puzs5Wlvkg5UUnULDPNd
e/nGIkz9BUspjyZtyr+vb+u6IWx/UO8E1IU1C7T7UopMBanTbdC/FXxHeqN2E3sf
QmkFZ9JVBhyIub86T5ncDF4868On7DOrddYZeE7wYSGP+gLfGryiCY9UyeK2ktLr
yqY3M1NzZOY0hB9vmZ5T/IoZJnnqxCvwM2VCvv52Dw7YYRT8kXtzKOHos7kZ3pJV
ji/9scusqu6LKwf5wjDeY8exbSUXwlSvaG2hTkYPKMLNhG/1HWVhNuYse4L7K8DW
x2gIIm3FYfac16wrrqHbkMcgE/S4aTDzGJ1o15Ix04odsmlt97BzQYwQ6+5s7TJt
+WQkTTfwQ9zde/ADDspwi4HFNpS1XnwsSXikstNBTrD2uPSvwu7o4TL+f9Coxrac
Lc3VDiE5jBLnm3mKF0LSxV1mF/gYXgWCuUmkDnWONlNyQBqIHswSuRqOEIIe3ax+
MSG9QT2jHg1Sxv/Hc2n/dpJwhuDH+wHkp8ZYfX1okJZ3Hv3rCyEgkgFMpJfIUVJ5
FozwzPE5ufA6/QdffOfeW+qs1S1hpXyaNub35A5Mn1Lifyl3KZM1R8YKdaGEkzaT
QbcHHkyX9x0rxfJLYS1dSEbqZBINEEgoS5FaXn8ozpO6FhMy+axVeqbmuEIF+sdU
PEKMJsyvqEue9o94aumxWx1e1UxHPioe3yOanPSwJBY0HhQdCz9Kim3jIVkN1q3C
JLA2GpTrBdDD+hrk6Q4ajsv9+uULK/VVHDGvM12jboUOOcZHsi5dgFVGiOuuJ8Q/
e+nNv9F7yU3ZIyMFRtPh5fBg5xnNEY9zlalWeZy9eEZ1rCDMOrPjxJnSwMirRxuE
XfzUg1MydJmXPhlNbFbNRmW1JdublxQBdxBazXGPHjY0GTRR28Nzp4Pd9MjvZ1o/
EhzdCq/zDgmuGc7Mw+tDoJRpMmhn+7iOkDuvHV2raOtU1cB5T1riUHZAnp3QvbsT
uMxt8DLpV5RMwkPFpUTrae5ATHNdSEiZVBUCh5rIy4+O20uUMCv9qLnnIGylXEmi
+U0N7vNeesHVxIw7xZL9+/qg6R1idwiyQkgwz4qDKtToaICelgO6LIcHRjs4KxXb
O0y2MhJvo0Q8nb3utFxeYwwGwFbrU0QEiEDAWwRjxN7jZqCCNNQ3j3jewYcqbFWT
P9Ys3ew3YwB0iieytnJeXhvisyhtPN2p+xCKFz9d5U+1wAjh1t5qjy7X/+3wXdVB
aJ2oHWzn2ZSQhulEShD/dhoSVrJZooNICc+010OCQcyIkZSn+PCz2Mio6NSEzAwl
HcxsUd7jAEucA1Qk9IdndjuRaodx+2Y18EmpU6JZzd02bVV6Bc3MQ8UsFFU1hku3
8IaDgxxz7Jh73NM8Sa56/4aByR6dX22oL1ildy4m1CBAHRjbNL/toLXnewrlg5yi
mVbnkvBrcJENMNyXr3xdgxgv4VHtDTYK6JSy3ecvJy5XT1TidpSF6n3K+ImdEoyn
gwAq5EgA8iJ43c3OWJ7Ymm1IalFjmPs4QtzEGoIsrzmqu4jdO0My/yp05uQswgDu
es5osunf1G2YzxweUNubv/XSpO8JrtBQtYlX3HQboeRaKz3Qa8yWIV7c4oAXYQdB
1Iay6w4dmKDMzzwgTMoc4sNGCb7cuBQG/KgpFrTt6BY2K7sw0e4jeugpRuaLZ25z
BM/0H3uYPfis0uTDgZOb610gkx3U8PJI6XHV1UdrDIqDpW3TJF3OJGtAKfWuak+E
GNrY1HkmuZE7rVTAGB+wfxauBnPXnFicMNFuegaDuMRb8R4EFcBFak8JqK3Z8Yyd
1+0dNyBcorV1lF8q/jB1M2BkoZIaqBs8dBGYiEF4gEsGfz0aKimnHKHDvDksRaUv
qu3D97FW9qPA9Gw9z/s5VX5PDodWv+CxFpEbhAvt2I0zq2ODjfHaDCGVyJtbH85v
PsX5r+6N8/BY9bsEhuZYQ3B+TMBrwHQdwiU5ro6NmnLiNpiOaekC9v8l1ed/fjWl
XQJAZuZ0Zp8Qm4Ruo6+JuZRwCCdfPn3O1ojfsaradVvUxpwqeYIG+Ax+fPv+lSpg
/YHXCJAwoP2HVJi72n3u/tui7Osl8Z3EEcU4/qqE9dQu0XyAtTwyKivpZqsE9OzQ
5CXjvMD09t/CrP8/xFr8QGsmgwQy5i9lkR38NEQpGHbJ8kKp/dhxeWckTrKXArdU
lELl8w8JCsepf9LcE5Tc8gAFdR9eyoUyzxiXK/Wk8UWW0tQJgKRuoccmMg1aUJ69
5PcEa+h7yIPPHEJ1ExkQatnbbqOPeYSEESwuUtHkmCFO2GEO6R9NOREmHS7EdiY1
bY5hjMrN+yeaHaH7tQdJeWV9VtjGQYs2A4IqY0yVxl4khihkW19hIKP7dtpyuRCQ
FDO9zCgvrodPNQjOFregLSgovNp0E62wM7k4JjU7JhMvlM9gCxc4dnU0zOqlsUN2
dOOGgnqn6TzuaBpqGcPtIWeAYwti6BWBfuiSlDCgc9x1jI2+CQvdNFyKhf2ci0up
C/FVRkXh6Cylqb4eNgafY9naHttSaNPoB8iUfxZvRv69WaGV5sFizVI0L4F6tKnZ
YTGm64Vn44PSZk8gic/lQEs8xNa/KaQXaeYar4SA0axyI2FD4FnR7b9OkBYhTBpO
w/kCS5ISEFVKmWUjxiZra0S0icvBSoJw0E8NMrHSGrkOnCx4eWgc1Qt+YBQc7niX
ty/e6NxCnwj7mnuCy1Hjt5qjSf1Ge0S0IluR8ow2XQaTu3mZ0X+SF9pH28r8aTl4
LkPcvSFueIOV8HaZ+Gqh0GXJRovAiB4Hvnf6tTfFLTQHl6xPH8oAyvtznZnHr8z9
ogBs576h8cvf98HGt0NAZgPHvd+3ByjYt1hmD1vWnyF7M41aN29P6Xi85kQCVVDC
DVtgxsUu9Bs0LRq6aHlR4dyGB7bkGmVP/g8+lIwwWveMhfu8y1twna5TmBk6Q8Xi
6MhETNDYjyP4z9YR0etDMd/PM+3NiMtU3YTq/hnCwuIERCNH8u2oEqMbGPJ3/48D
tz4vx21TcNCTK+DUfryHqIt1HgNAOc9x+GqdMgkpmXC9zORBPIgG8u9Gb2V9fRQS
Sv/+U044CcQgmaDUpKagkPodoJUub4dkMLToMKxp35obVmH8lcvT8q16Bqfetrfr
oJ3exyWJV+fHrsrgedIwghDc9aQtsIpFy4PsNvc3DGx4vGb9ZD1koGQ4nHtwyKOn
pnbNMkoN936Ps68JlNauiP1mOzqzjh+YE8e8WRfDdaAP3yagNNRixtg5j7W/Rv+f
JhUxHu4ulV6HEtXVPq7t/E1/kAVBOCX/s6JGyqRn4XrKO3C1/Ow/0gnX+1Ll3hIw
nK+0zenHKEwm1HFdcg9bqtJAsZvgo6NdYUAwqmQpU82T7n5NgtfBh+YdPH5ApQcc
mawJikBBeoI8798Nc6itxBLQKJNt42dtQ0bycOiS3iiTLX9od7C1TXQhAusaM/rW
T/6d7iN4msrndBi69DY48lrPnzBf/26NTeEB5UpYxP08dsV43NtMN+PN+YwDZFES
PSgwtL+W/jp6apB+IMOUQqh4Ib9RQ5XOoVxEgtVWCw0Xe6pAhr9ExceX4ISBvhT+
/E7g7h/PQNevkqQDlWx9SmgFG8A/F75ppVmf7BOThMR1iciu5yqYtLyJV/QkT8la
AxOA3eOqZUd2iy4pYF1t76D8dT+GtwJWobX9XbPweZ7lhsYRRHJRqCHjtHvlT9dw
d/LEeuqq0fJFPsdN9hjtEycN/8T/jrnP/6FEcZuZT4fD3qR+QrfUWjmvYW6GBwyR
WxoZEUPi0WFNIX6UHAoCHSaX76EForszGYRaKVnDYzBD1JCIkItSyj8V/yEuSuXK
HrWMLV1e+r7ejhujutO9YNXFmie+pM2HSJO44f9n9xbmUfC3saLQR72VKpC9RRLl
A3TChfzYTIPjKv0VK1fGrClMge3/TGwb8I1p2N5tLMpNZv0XRSpJM1PVC1c6i2e4
ehKNHi9U8u5yD0PpR9LK9OYBSAnSJpzKn8O144BJjuolf3YZnn5rizDZoTE+vgXJ
wh+pKUJWuimpiDzVqRAE6HRcojCRdYiujtotzMyIoG5r+ArfGHLE0hHpBLOYWms5
XdZrO46tgmDtlb6G66zqFdhJ75CIie+8wczqmkpMr5r/iGVKSDrvVdoj9S8yL3zY
IycT96Z0pFDTc0v0M6aD+9mOSyPk/VDBOyYMc9r+JY+SpxIBGj1iYoZR3qETTXuV
spK0wDI5GH6OglCX+KSAN6ELVQ2Q3cJMJru9UuTGh27In7zOXJn51BkaaAJsP/8j
mOQZcp76Ic99W5WVZeAJwQWzsirdXEFY/1pgBHyb6mViVoasJ9KXMGgxEMDF6DmG
EGlmNPoVzNCDqzikfFcuJLDHCHVwDrXMeUf7K9tAAzAQzO+BhaWholidOS0yVech
HYsKhiJdiMvRLDtN5avgyLV3sQCFjqkQFb2+BKQK5Jzdmk3dh5OTRQMO52jUCtHl
dJipy4Zfe8Nua0OM+4Ob5KOo1X0jgPY/2cb5h1mYuTYSoxw9LU49IxFg0HBR/044
9jidub8l+aaeoQCrvhYG3WR4LaYtzUz+jHoEKjnSyeor1AS0oMUSyFPYePNAJDUr
UIoTXnCiSzs380XPeFOswWbqbrZVVkxa4MIQj0IOXIn3rwO+//9sCB22bJCyBjLk
/aztKV4FkX16mYubLFC+Q2wJ05om5km/Q1a6xI2VGj/T7qhUq+wEoex+PD61ZQm3
wl+i7rIIv9Jy3cI3aRgKFU7LnHServ8jhOpjrrvd3LUQnxaa1y9LslNH9vy7BPjC
ts+kdEimT4HS2KAtprgGf09EK30VOTq0mwYNwjOcSMlJNu/tQDgSvqEc406SJbR1
V7eFaxND2EZ8k74EmvwQHtsvb0/pL3fbLLbntDTWKS/v/+RSgacwc73FzV43P4Qh
DxzIpcFpxdxeIpvu2HTi2i8hW4N+QihEZCkxV6Vxecwn+Me/r12lhgkUekFVCxyo
65gsym1IIKKdXWAtGzsfIP4x1439jyedpIOcjZAxRVRUi5AJzLeAqYUbwhZPnNiF
BnyPesnpGsBpvK7Jut6MNPDr+Xikqnai/jWfLRwCgOsZ2U09P5nAN9nLlqqX9wIS
fH7jAF3Kast2yPFI6ERmuLEaB9EQ9kHVG48xYQdAoP5uzXeYE+lKR4BaLjyDIyBV
Ll03zYsZnc/S/bRGryCFCDRmFJJAjKqULeeLdlucWH93DwnqECmhWBaR0ge4pPEi
KRFeosRjrVIb4FsaLyfN/50SHA7RHF7BixNTewhZRCGoSIo7nw7VhKFFZt/2cozX
FU4gv0EkwrKPPPG81JcaY/hyU1ZZScQ8bpvKnEjP2sFkAWx9aK/nSx5bcuNSW8D6
bvMNkATehPG9v0TrpixMv0H4fjrnPsh0/XfAAINgIgYQv18SQR7eAz8Zl11Sv8uv
WegdHH3Sx9tCG9ZDd+vqvKEg5Tp/tNlfqAtLr8WPu0fCgxJLk94yhdAUtYbiLQRw
yzyVvFEZYNGx7/KnRDTAKom3HsesHHK/0a4z40UeMiPexsfxeZmTrnOtCBhE98gJ
W3VqS8uQFpHBBR0YOxx1sGIgtad0qFj90NN2x21CI07oMG9veaWK48c2gEhkama0
+roa23c0Vh4fwiBhGeuVZkZRzCCFra0Gvx7sLh1wt4m64IiDQJpigEuwKHOnsTwr
arS9rIxYjcpMgqzni7W7+AItBvhNYV7ey5+dye8Rsy4yD5kVIEHje0n6fiIiUZoe
wrr3VyT6uG+iGQrv2MAgfVhBCv5v3tspRv1ePC95s2bvs3+xCx8c/hzdhO4VVn7G
Xov6k6/VYIIhUXjFiFeAxm/YZ00YPr2CAbbgTfDsJ2bUGpxtxIJ7h5jntoXFjV6G
yzInL+sLaIP98VLUxPhRpkSUh3V2I80JTFeasSnApWYcs5B3GBrlQYCe7VS9vG9V
dDZMxwgGTiF12OS/+94PcxgkSNW9NR7wE9wNZDaWzs5yYfEC6alv7L7ycxCXwy9h
tlwgLw7pi4H7ZaE65h/BGZBXxKWiDxVcwzGL5DbuuwqpjX7hggMjx19z6AgloCFu
uzmbXNspOnH6omkzqjRcWmu/Xm33Rwr98zpjNC4lWtOgZjUjbGjVkX2HbIPD26bC
uqjB7VwoW5P0R5hlneKDv9KYd3TPOG8A0RCH5ncw97sz7laAbCKudGgAcBeAPZZa
Z3MXnkZlDyEvUDL0FySMRqPftuSs39r2agI8GQRVOUxRT1nmECRt1YnmxJDoTKlj
kTptFcz5kvr5aCFehBSIVjopFAJ4NaMYCtD+SFXYvrnhPftQpvKh0m/fAj6jsGMS
zBCTz8lQ28QSTyEMxNzxKbC3HFz8rcnrXV7QgpeeaDT18vxzAie8rJlY00D8SFKa
0s9DjRWOrFxS/lE7a+cO5f5T1kB1u2vdkPnj6XUnyp56X/71zvsijX6hoinci0uJ
Ps4vkuzNFSFE8L6vRmRxJnUZ12bVW7IVlP9ftV+KGi9ydCwTbztWse5Rd6vOJaoG
dow4tjD4kPraYiucUHIhgpE2MtRgPnvaffvellDX4WdArPCjiF1LToKV9YcZ9P22
CwauN4SbCRPRQSX027zoVBZ02PwaUQK0DDYGRhga8u73QXabC90OBU3VKtYw2ZaQ
V2S630pwjGm2eoi8t/VkQ18zvizUeHLxFt2ShLRbAqecV87CB894WlUpsK+m6+Rc
r3HENfU0uvP9W/Xd4wT0uv1/1yo/7k6YohwlWtjhUpXG1qxMqh1cDufu85U4QvgP
cbITC4tskRSn0LhL5DBVA8+ctSsfSozhgEnR0wIf2VulbLNUNKQmC8Mm5FnDgGEq
QTgLz3KD5OxQqnj9qBJAX0/vChTqLMApJD1pHRQrMh4K8zIva0fnFGPC/8/e0Q5e
0j/e3woixxQxuD2q8zUarNxCRBsDtGbxUziCag3XP9kQYXU4VrqnOh/Klq2uduZ5
iuUCVRyfftFm5NfoH9bfrtGEnKGut7IIXwrUyVCzXscX+MMTucEO2zRG1IjMxkWR
opU5UgbEJA8MkbPkMvCAcAtSrwYD0XD4M/C23BwQQY0M1ao8dth1KmiM6mHLrBCd
FcVHKp40/KqPYd+EhJky0EF/syLiR6uq2TlbOcABbbm0VxuORA9PlSX11YLZRIfF
X1e+UXVhGMHu+0cRN0iygQf1xDrY32/ynoY3cxtpm74BCWUbDuH2MPrkgGBhClcO
LuKfDbkaFKkugVKraKaDEJz+HYYoJhWcTvmYHx0syHdD8Ik/+r1UvqZu0as4eS2A
ZmjkOO7hqLK7suCpAsmVEAxWjlxjHVpodyhrH5cmSJXRThrb4k4yJZF8zXfPmDBt
gy/apASkigYsbaGd9fD8TF43PVmASnPj7rFjpNu7vHIQ8XQC8KGegTfiH9DpFuhs
tacW1XD5iX8XEtOiYccBoZnfr8v71T0v9fCT6b9N7AnnllRaIaJEq9ZmMbvkaNyG
9t2osmlQkw/ohCrbpvGfkC0G4+iup7pw4B7kbWYVELhbTtg3I+NT6sa6LFAa5ZA/
Z1TyLqIWxBgpaOysLW5yt1a0tYooHI0hqw0ZhVfCaL+tuSueAtq7GmnI0LIDXszh
bSMpXChNxT4OABJwaHK25CjTt5ucYGyRIBs5Zn96jxzgpqdkNFawsxPO9GNGSE4P
UuEb1Pa35z09YY12SUkL3kfG9+E0rtaOQpaDmsZrgn2AwGvYxtbIUW2KEnHqxAIa
dR+YCQ/U6Zx6mIiTqEq3ZJYFZHABhceHCZSRcmvryt2GujTAzu6zsTwqkqQJ5Mn9
l/q9Lw+g0TXR2Wh/qZWR0yxXOrggwQabyA7Z8x3u2Ix2bb6Jt+spC4b/CDOBqfeg
04L8cd+IvBnXNU6N0zW+0/ZwDzTTXV5V2hta4xcdl9S8g4SQPfSECm4V41D1gRXa
Hu7w7Eweiff0lGD7BiGGYy9CGxN3KK4+d8aLcCFf0+MdEe0q/9aTkM9YEjEJ8KkO
efcVRsG2HHh2gxHamSkvUVAKf+QpHNfmMCUonAdMDUCLkN26WPJXcV2AGmz9Sqr7
1HXs6AR3AAIzd8qRNCkcae0/21aZYJizNNoBuK0LzYcqVf3HjMslFJRm/xTo/kBn
Ip7zqgmlmzbYWrwTpKzxkjbfAODAplIML+nTIee5NQ39ZwjkXJS+daSIIesG9m7Q
lvsYcpZia3iShWL6jfpD4Sffc+YyvmEeykuO0PuIywnXXD7dU48DGA25vsaPeoH0
dZizPYU1aHIHlQRebd2V2WM6dZObJwdpCVmv3nL99ovMuzFzKQ71LbtJDl/tF2Y+
NKCV5han2nBBfdCFqrXhGj06qcqXFU0Xo4QjpmkBDHqRxDlTKjIy1KYlAgLlu04x
QW+WS2MkI1qLkqdQe/NronYFi6N68OAAbteYxPAT9wdCbyBCBUwyDcb7Dt0SZk5k
Q56LqJNUr0cUo8xT6F7n76iPV8ELvJ57+JtM0VTYTQO0uqvp4/xfzqXxX+jqGGwA
Vk7u6jIrrikfgPIxwmJbiteZ1Ya/5fmTXg5A+ye5sTmAAOibHEiYwH0LZmWKRbPD
GKnC15gm067Y4FJo7rdL37mieYkPLEQTeME0AlEW/eeOE7nbrhgn6eF+LJGzfhQV
Csw2/bzm6zNOzbI/ZnxA9rVRTGXXvb0FRBjvonz7mvwJQhderv70R4Pd8OOamNbF
N07a97vEjs5X+248z+NFjJvEcApB68DfJa0bS2/BuWM8T+ODJ2FG79S4TC4F/kBB
bOZGd1TdhA1N2QpxuVk++7MQKgQV67EB+oLURRKIPSTyKlzWEZB6SDXkOIFxHRz7
zU2ozOPVkVI0j1s+LJ0OAz9RaymjPuepzzZ7jTDuUBSxRSAmqR0M7knCi7qGy4PC
TzdiGtLi6fvvAH+DGmPzt7F6MyepCaXhETWKjs3reQzMpx2bf/e1Uoy5S0voXH2U
jLoyyrIQndClcs/oSZ3hGwWxrAGmch30dGjkRc4/rmO1YQqngZ8++RV10npC1l/W
L7bvJrRIzpqGSuNME2UTPuxY1BmIfe8SazEP/P8cDePxoWxa3L8vUbwORRBvozes
LtZ/IoJDxvW7trSrjt4GbWkiDiX5GPKiCbKeZQnGpf6Pnsg95+ADYbef202RxNP6
qZci1nVFqjhLl4qVCZ6cj4Ov1QEe1vw7Fy/blTx+HZ6WzCR1NegGmw6lmzMNKJMI
LsP3pyJuP6aXf5Ip8rKQbsRrJ1uZchng0maD4tuotQ5jCjT7iEMWgMjtisLXW25t
d6Bd935TSq5IXAWY5tcR4zSIYuD2FZsXzzHwah9HegbUkHKWJ3ATlNSd/1VVtaMf
xuqIU8Q7fi7qVvSbL767Vog+PG1dnSBU8I8jNYqZm2leWxRIRa8KoTr/7gCYyMW2
L8D2/aaB7nyZmjd7ov7w0MExC7O0dHjgZ/9v3oAUeSeV/+0i78opAujoM4uPruWE
nqPY5aAgomD+0MbB/hkq1AB0tAA0zpt/zT/hugJV3F9QRip+knsloS0ovYp1p3aP
geA8YBicEIim4Xa/XhbBMqS36aJDEXPaO91vNDrI4Hrqkv5IKXJOHmbTtrWaegBS
En5LG9Sm3z32KVK+RUTxgUJJsZe7f2bscv+AZwIPNoZcfbq1IH8nF/AXXLZiZSjP
Zd0T4HByh5e90BhKvS7MqLiNObDAo8UxUeQ7+QDl6H517Hj8BaqgJeaHFBaZ+XJG
3DMZKICDCWeY8WglU1awiXJ0/NL0HwMy+T2VGlWXqnssuJlbofIx/urH7iZXDILp
YMONwMEAqu71qKQBE61OjPZ1AXr2LBfFdAYXXTqbK0dcY+lk2Wd9VXR9TyCchfP5
+vBOuqZgfyEGQtRq5tcPRWJ0xXncLX91yjHVBfI6Lpy1InJXLULyEGW05U7rBeor
eGK77SJmAe5FlsQ1UzWMFwZ/TRhMOEeZVca5qBEr2DqssgjvBiZIshNwf783/00C
5XAhEcECqDyss4kpj9UDOQ6ybGEpJTcbLtQMLiEeBXcyOV8Lrhs9+JYla0tlnbGZ
dLc1JRuaEroWlucojUYbaez3MXrr/4cNpzjWlZ1wrdGA5pyp1NzjYz1PqVMaZ544
N+BEP28rdcbp7nijVkQkOyLDsgOVwuMaZDCDQdUX2BbkUpDl4Lz/iAWZyTKUfn5M
hMKVlsdxZYv5lxVZMAZdQ20Q4lBc51Yma5Pb0j4+6LJoQAAcbiTWEKS9oyhaTwOm
WEoatvg/kUUG+hrrQ+9E0gIp7l1xShQ+otVgx13AqAXen9aV0H6KD+LkDTxhWNmO
KE/c7vQbQW4pLT8wh/ezIG11J9mgFI5oUmtz2qGN5xfvEtj7jaKiRip1+wFhkUMG
rOY3wQZWOnkg+m5Pd0YXrt1aYFooDNMLWQgjmITo+2bDK0tEO1u7cpJd988kGtXx
11UITG/DKLoAo5imUksAVfKYyA4gK0a1jpLrqJun2RacTSjy19qN7uV3jJ27Fehb
NyYlmJZq1OJWF0f7ERBdFV3EXtY6lw9kwbReNhlmp4QHpXI+gXvuocJVTJlYUWE7
eHT2b7POiJMsMUMKV1bu9ErKhMCkk5yXQSZ2ozzhVqJVPSZZ2VOYZ52cA+rb3BcE
JQcsXgOqrvAISHg8P1dTkpjEIvqSQWaxMUN++yRACGlOr6X/3YEKfHWfX/oo7HHF
SbeOw8XtEntp9+/+qbKsomL2riuam3h94yY6nsrIi+ri0Zmj/+FGK65xp5gA+loQ
wzSzoJq8KVTfIP7glkVkVL/GylWIb8GJFVYodswktnM8f4lF9y2qwpBUxHmIgv90
1aBVgHWxPJ7H9d2+RbM8EgT2Tg31F/6L/9XQu54y4rJURdMh8sH56Sh6VaY+UbsX
JhdNXcG11Y1psS3xd3trfF1tPhUsQPGJMauwK5E8cbtBKYV8xh4ZJCcFyADrR6XQ
Lj0VCzrwH355yOaWMNw2/RsCKYFVH3eN9+RAxjlUVrP09ZvdqzpYLRiEVOncll3m
jysNFAOaZz+TC5gnBi1dBIkEgdgnuu8bDOQd31yN9hOHRhf+hKbHod8kTtWUMKzB
t+9pqMtOqfVMXWBzlKa7VN7avkwT+HjFL2UX4IgkmnOMCLcWmkaCS3STpUHOKnGo
j6pJA7iRLWXQCeu8KiIwOrHMMpvQ4y0auybn7vGVjKhEKVjpOJJcSDnToNxPNSim
eNYC1MYaHdLVm1luAfOo9BZSE09FrY2ZNh0uSYFQKqeibpL8mSSzH6wEH/nD4nxM
7x1T/f2W5UjoDNKSJnlx97M7Oip+yRpXPjUIvv62Z3DydQ+Mag0Ec9JlSaAyCh9s
CMGjMkY9duWrJMex2pIxQspptwGG2nsWljFbUgRWLoI1HXy1AHNcS3UvXCF39jc1
eoLKld0ZSnWPuhbXcfrJV9kDUhxiyMZA982rbNe4skBigPWHy4oeRxsoF7AvuEWw
1zRKzBkpb5lu3bHVUfhaxCxJNqa1rCAvFZCtQPz1k6r/fyvuy0RBLJSrEfGUsFJR
Z2BukVsyzFohJLUD5deQcBopZD9+g72ueWhRIkEULDx22DI7+4OSSbc4MdS1ppFc
hts+lEnt5pFhKMcK7cs6e0poXAqwnKKbFeZWNBwFuXGOWrAdo7T2T63XngE/B1MR
bTX75zG4vtCYJSawNIHdyzvX2sH4F2GbU09YlGdZmW4QuZe45I3QDRi9F5VtFvIM
zXTQvqfZUu6HJYQ+2cTo+WTEmquakQcqgRJOZnm6j6an7coyc2JrCn2VP8RaDHMJ
mH7djRM1yKnyS/hqWiskvnd+XPDIZjZX1/D6RgZpLNCzyn9CCN/rl2PtUBsGartj
yL4Zy62f3ndJGdwI7pmyVFbzUraVYONoyjPMOCSmOq+c0/KZevOPiuZtDm8pBuOr
8wUtKnI3MVyoVYFEGtq7jZzciGRhY8BCUG8CjbOuyUn8Ssh0kt5Y7NaOvPdjF2VQ
2gitD9RVMagJD0e2UsgFPVTba0cocvIn2DIfxluMNFuvNYcIpNZafNWIhc8fyQwm
cbULLHWJBXiHTO9/tkkUhddZ75HZHbXMZHVoP0rhyVAlIMm1OPhUgoUTFVO78HSb
zhOuyy5r1+Y1gx/f8C89QaOWkKzxlOymRHLmQXijdCJ146f7AGN/UGmODvciuh1h
7l3hzb3MBFZOumGBwQPArCQlbe6KuQL6dfdYfYzUGWsALYy97m7OH1RdYDLHS8Tt
TQl71FMwvyzkMPFqpq+LclzovagJ39QlfkQbfzUHFjzuvD18NIWM/xEqTH5JJrqX
Bk/5lk1x+XC2nC+E+EfUKEjnmP2n1InWcJ3XByYGs2P46MQT/ev6OXoOqo9eRg2g
b5PRtzgKTCo45vy8W5+ByjpgjpnlM+8XYj+h6cdJYn3YCaqSrqLMX/isY0VxWNVb
p7GgPlStGR0wIntV9OMdNxB7JtO9nQBtNNa8f2AiOHPDya1AjsZzZSFQPqN9r30U
dl0wkH/EmUkbr3Ex103kPzGkVmf7AaBDlVChBh1eXdErSinWOukjoj5sb9Bsf1I3
Ow9/PSVnKBa1W+LE6bBW88Cux2c6nO19WOB+nwLTzlRgnRwAm1yPscTPgHtIsYx9
ycbvMewjlzr6ZYyaMSBpk/dTh6OYnZgVzq1b175czWgCAxiA/2DyI3zf8nR0Mg7u
rBFNANbp9xjaw9v4fv9FptNAnWMKYB/DWCINpq8xeCEgkl9I8j6fWCeVvYMDuLFj
DYLbJUuIJlIXLYuwuxWT6HBJG1/pclGZy0K5VFmKdsFYF5VcpeTAIoGMPXw7Wtp7
o5KF0IsJeT0n3Rv3F6z2otyTxRLL4XKPE2PUUcJDF2X/qiuSamijfWxMXxEecJJP
eWfCHGBdTc279UE7CXNilQSMlYiKfzNHoIR3ShWjVZtgzyn6oB70KkwxNVvhLnYZ
euBAoLiV1fhQRpPEoqRpAW0DYQZR00zW5bbOqhxeqKlf0+pDQhVvAs0RqAoSBWc0
xPtsieNHvwI5JWXVqfsihc989j0JPyAf8m1PLgM8nX+5Z8aRcvzgWb8zYKwLnZTc
vunKANpIS8ki4649DMEfNmhIpQ6Xyob67ml0NCEficu5q4ZsQ7iWeirsAKkco4Vf
jtu8WnmaLP9zjSNsnhqK3uzGAxqmoEGHT7+6F8Xj9t/h/xKHXpZWhF9dP9Eh00vB
4Zw0xXPG8WCgQFY4hOgoA5EAPSM6uM/uI6iHBRSELID9BI1c9JolCMBjQj+eZQJx
6V691fkbag5Tt8LXP6lMeGAz7MFfEiyKHFp5rB6vdy7H3EmPF5yLIQvXwv/ziRR7
rZnmTDjzq8krVKWzWDervz9uSmUblsLZI4Nj1JZclhaMbinJHL1P4510Js6t/ljJ
P272abteMIWJX0IGRolv/VXAjCRgT2Yo4D5j5gnXVoSzvPcJTbqCH7LEWgi2/fTe
7058+6MqsNE1zX6uJglppjn8XzbBdX8l6iy6ha7PBDdubMY9Lx5HcjTk/8XKjlG0
1uPltIDU4bv/+p9/60f3AfZ+uNjbbOLcquA9C1ASm6gmKYiMzZi5or3p69628MV/
2OkVPEmBWEXvPUuQUtsPL1+4l82cR4MBJ6NVlIci3ZDAgDSJO/T8yczqfD7oi3vu
zsyFDmG1jrF8hGabzH+/GtTrLNnyms4BqUJj7R1nsd+KHHwROYfYv9xKLAlAdK8c
dwRQLV9Fgcczr6uOd139Ue46VFWLmq1yoOoV5uGoJZ0WkqHUCC58SiKqP4oWWAZo
U8m/P9scyOc1vh3cvFvrle/Bh0iB7wkvegbDB74WZcrmgiI9yZWhR4ORJzdrk/y2
OJGyI26RgavT/Gv/piuwC8u1X3iyBZlGqb0bm1BKI8s/BR1KYo/dvEHD0m3V+Q0M
YyUAJPmPIfT0Jz9Z8V0HqAKRrMJxuRTSKSUf7D2DTp9rJ3BASSDBGBGThQ8NLxL9
awoT0wFAjkMqVhGTiPkCZeIbDeoQ9oNyUYYnXsnAOcDuxw4M4qcOpiWaQ8AdDsmr
2UIdRjV9p/GNkkgX7T0wE87IVCKQgaLSGWAhWW1wr4Wm26llPD/LcqYvnbvVWUxp
16QkHqojKXl35uzd1MBnGcZ4PFrFNY0vTwTrNfP1ApjR04w3Se1XRi4hMaKd7lIk
8w3I/Z9dVC3keenvDIM3xeF6xGFZKoZThcItfz7OT7LZtHeABpcPSIYruhPomMGg
5eF1RPz4Q9UBdLedUMaKi9t7TGLTQCMI7m5WO7VMFjGMPCWx9X5UipyxRlDMQvP3
gRebk43njx2af0lWXJWpq606Gc0240mZmus7uTHuLh+lWhpeJNIaReD793TgvSmR
P5jXxmEg6fYUdMaEC6dVnqIhPHx9NRoK8STMUsLdk8GA3E26MJt5Xk4lvvC+e9oZ
vM1E+xPn6jJYuGnsgvjJCBVMlhzExTRopTZNex/2lk5R0kePKr752R2jg7XVfiXc
sbOtsm/xcDaB25G5RvxAYds9YBWwaDSoluq5na5lhPXIgyZUEUyJPAvqsMc1nuqC
FG+fGZ4YJY50GUgNlxIN7ikTsnAYDyttzd1vS371Uxv+W9NAZnevVgbAjmT05TPl
W4f47He81wSYOjhrBEAx5u6ao4yzjWHYoMV/DAqhaYWkIVoL4gsRVVnoxAIXu8zJ
dmyG2SHG871rMB8oRTeqmYuo0gGgW3RDDRWhlT6zLwEjy/UzUlJ6gLELz+U7O/C/
REEB19t9T8aextNZ65Xqi8IRo2CQRK5aeRJDkxByI/hvpLePje5VwtPoXt3FmOju
IGHiAlqiczA7b+2e0QXqWmq+/64f9nRppaLr30x/QiiGkP60O5OfirQLO8jzv4BW
/DKGFeDZUoNCgvSa1rPqeBUtfA0un9tImLRr5fP5AV8U7Rht9ZYO9qiUtDx/ylOn
mhEMfzpq7ryxGHX11LEF1sI+Hw7kO/+4XUaDdgAed6je16heNBg0Zb8e1q69cM1x
k3Y/zN6M1NFGUb3c74f7iuSQE9YHgYbnylcoypTkEJUZU/6lDDiXq4TiYmYRwIBq
4qm+6PhhK9Y8SPUYY48juzTjXW61EeIQx/uj88yAyfUxi01NxbpNk6+j/qfbEIE/
qLVvVFhSXDp7E9Hkiy9y2/+GbapSbE55E2cx5Zq333I4A21yTA8MItzQpsQbDA5P
FeElATudpL0gsawzhPBfHXplrQo33AaZc5suZ0/Az0eIyI3qQLuvU2k+bGvH2YhN
2yzTtybnmW1wW6yYVhrgIXqvdErwZW58EzzrcH5/OCH5xH0SaCWOxWfnUsv0nU/q
7YsyZZ6nNgHwShKPXOTnSc4NG3pw5HaOifnQ8S+WJuThCjwV08r8AYx7uUxrxgLE
c3YvkZUJbnW78+3yD9x83sWsvWGAiH6tBtq5v4DrHGW70nOPGRsGisH7gc+8l7Wu
c/peRmSh8c28E4yZtddMnwXVmYU2xXLbmGX14KIYOYy9QZNRpDieqzXXDklZqGty
QuDbdSlwLv+ZuIZUA4Oz0TfQixlIvnpR78P3KdnKivRP6MhQs9NSP0bkQq+qW4Us
+vpdqzKJT8mcO/5eAUsEWsvDAYCNddWZ2NZpDVm3d79QU2F8yDr2hHYksH5I1YT6
/BO8geQ6NUcp6vNDCeZdLJ2cqGp5+Iv4n7OnzBxZcm8+xKRv90kSZfcq7wcau9na
6bHjZXKdXl7U7F8gLuchUGddHQTEO60ZJ9Sf0pGME25+T7STmsFygHYLLt1HNZZ/
9RViVrYmXefdEBUPkNWEig0HcLmu+OuTh8eEI0RK1TBM0EtgOzHZd+hNMrhRoGRB
OA7MpxBiYDepdvg0a+gWWE6SjN/BHKt0yiJ22k3j9R7rz2995UdTZGcJnNIfPqT+
XBXTeb+0XY/yFYQUfSxd26YuR5qmUfhNqTA6vkqFqjhx6ihYYmTowJLNc5vuSAaD
bdg/EFt7ildeLxF4HwMwdDqx7phjQUabs6Uj5RPUruojvjz7JaawmtWpxQde3ysI
4dpORSVzdcXktv6aQk+mN5wFpJEuCzFV/ChfyqYxrl+SYTrk2EJC2LcwK83noHcu
4nwjhdvn11tt5vT5A40Vss/pdKzxckr844Ai20KjrxcygbqyZ3tYnXMtZgIaKiyq
AQH2Kgw0MvfrOM5KC0huWEEXFX2x28YL2xkdh2U6TdvZvSzBndF/vlNEUyxvqSqD
hO8KljhKv6fT385WQ1p5SXUDkK1J7PsD/w01mzOUoZWak7jAsaA0sy+XAJYg3V92
9z6XxK9Qedkr/xlQrKrOJscG1OD4msBJxzndZjkEeEniD6McS2c3qo/ThOWbPBTY
mC2UsJ4qgV0AxZ9bPeW6ThYe23QDtjMh9oXNJDSsCNkbpalcwGLGvjsaEC8HumoQ
6dtKZ2PJ9sDr5MaQaUC9OjhPeFH4Cjoq312VkHN+K4IQVERQCNdgWHNuyyYsFx4Y
0ozAteKC4ZLcbNgZ0/aQL7DtYmAOF2kCtPKIcVtLj5hfYHvSK8PXGH5LFN2LALje
yp38Tfy216T2DoTwPiD7brR/3z9dT1ARvTsl7K3J3HyUDYD6ftkHJdZHd3KY9R/8
aht7+Zyji4J5JDztk97fdkV1waoZggcqZRQY1swMdknKPmUcxiqyE/86PiCWLiKX
gz2nN+iz66/10DlF2UmyCqLEVdzKRxuNaR52IceJJ8Ah7q4om3l6ktEe8ez4ZBKX
qZfOHH3vrTH4oYRSpZBS0yKy0Q5dQY1tJOSEKdrwERhfuLmwwj8yk6rZFtckWnbG
YMbvNdY37zLp4uljuGwGbTkgeU9cNb79JsSmqbEflWoLgEG5N+v0iEnvgGMkzm4e
fcTI+Ana6En0djyomr7kaD0nKPoVTqOIlzfX+xgTgJjO39l1YKQIDxaSscm3ZRQD
dGDEWwjTNKs8Z1Q2a0TB+UIaP8PCFGaVafJdRc1tn6K5gEKKi2wuRd97eGk4ag6X
8xjsNjVLO4VAOg5PxnewFCCfnss9tO1yVHRExA5KDzMTq1MdKn/qqfE8Qqe/Y87q
Y48rlOTdYm0zRJK+K3E0aIk2218AeaWs4JCS4MLBarY+nEgCGg7pY3ScN69gD8QU
igcDDEibjciaFuWaqPmE/wpiQpNccAzwh1YgNXp7Z4cvMrOXG1r5hpvsg73ifpiS
2FIz2jAEuR4J60DPAm8cIBFC22pqD5fAEedQoQTQ84OsTBU7IhHApa73/gHY4gHY
W9fe6eZSw80vPoXr0YeJ+P9GSKyq+Oha4sXtLld+9p/JWaWjmX/YFu6hCtvdo/38
GZTFNgGByeJoFmimII31z3FxodIU4XW/s43wljOilJvh6vQteJAAG+5CPm03G5mK
shgdsYa8mYt6cdC6JB2wKej5r2Ia3XhzuBrj0/Ex3ZR5bNEY/f+u+68Y4xWKTPy3
47QrG+jpR/xB2jXNF6KWN6axyu9B52gUBXCPnF4A6iRRXWygB4kxNRVLL9R0+c+U
CJXDEugJrdambcWkflKwpK1ugc7bkOrE51dX4Ip7rlWgLLgdl7pasoOATpOdsnW8
vEv/EyCMXsOZDm2jtlzjNiKA60VJJD1RhfNCLBe5uW7B358Ox4Ty7XU39agHgMq+
QEzhjz5bFx8JqjcHDn9KsgVgmsUnsxMmWuBg1PU3oXVOsu99dR1ZG8YDLJpjAHKo
tc3q0L6EyDxzjKGSz9A67xEczBU0iLNQfjVgVB+/OKSmt59uPY+QC9Q61pANdlgy
Op3GdZBDpPdQZ+O9WExf1rVSSQE4jwrIpMyiv4UnR4TOP54z7vLQ50W4tiY7fCgb
aJhy+CUzLOtu37lOMBeaMDU1BxIli0pJKikBjni/tiJhm0yY35LyKcF8IIbPtlCN
d/Ylv1gyj05k4PoEJj6fzkjpSjsRomjszXq3bilogVJst9Sf+C6BW0InvsW2nSVc
APJB1Rb3fgwrPiLiwP0uYXfAf6sQzGa/p2ctK5qCzTM9VS9A48GIPz4+I1xN40Wk
dChES4aFFjs8aCrPS1GvnTAX6sUAbIZBkJR/UVBS1liyNaE4RHBsPtOwYtm4xtQg
wZvzPZPobuG3uD2c4XOSM/QyqrKJ0npYzNUhrQxMNLGbisJmxYGuG5u1zAX/c13k
sIBTgP7wrvDeXT80oZ2k7+sQiAGMXQRroc6JxS34XKYfm63AmRC1uNg47RmYE/M1
YaDzZGpe265nRocjFcVQEJCjJSLkQZW+zo2KtaHIMrqbng1Pf+dufbOwsnHdEBzC
1baKl9C93RsSIYI7eQrMt90QJqih7KxJqncvNv7dAl0mZOs4wfW9/32nb5qUBXUL
ps5cpLOEpNOOLSP2uVCzgERfn7xEAwjtGPpnig50GcFaRnMO1ayauxf59EpEwdED
iAd2SdaEXyHwO2lQ8QsraV2S96ZjWZvG7SwJ9yTc0ZeYo2sGhvxJPi6QEqczV7cK
xrNbo/VzZbRbHTnCGp8gktWb55UdVRqbcrm8WYKFBq8bSksAvcCFFvV9WEq9YOgf
l+q7r5pkh2Y09Ikb/G5nleVLnH81mEvXaoLL8QX+Zvz9lzWfullqsE2HONmPYk93
4RzR1xThFFXPtk0sdVw8VWv7uggciKGs4TiI3Q+5R/giic3ABeq1H2LxKtHn79RZ
jrvKrwG5WiXcC3Cue1gXSP22z80Si4wsgspUDsm3sKnAAh+jRWYxL7qGAjT+npdo
FEWkFd8zdRRjabIfhAD/6Dx1FatbLolbxRyPoxcGx73mjCUFxFsO+TwF1AvBEAmq
abL1j6Mzq+X8aqL9Os+/pKt6AfDEvcQNMJji1zK6LJVOwZ1HO82fa/hdwmHt9q6K
VNHMApwS72eJv6BKwcooUW3ITooL9rLbvfzLXlw1Nx+D6tSzXRt5xnc4bYFgiIpY
XGldEQIgR1wZWnK5xXHsuxOLqq7Up9fD6PCyEL0l0ccfPgPM18pVqh5A9qFN2z6N
E1DXCMOlofyMw+9Db+F6vIPh7C6to64EZf3NsNRtNmdIOb+7MjS+pjAszF2xlNnf
od2nuuzrTSIFnkfBvIcfOarOWB9dlYBkJvCYYY4IGzD5naBWQ6c0fwzgDi3n7vrV
usOxT+UFZ/F+XUc8YPcRJ7E+7gOCC+2Ty4/8uXjPPyfUlKtCBWFZ5HC4mvUbB2bR
pxAWcCzLK/8R93wP31NNuKNVpyQjEEI+eZSz3gzBxH0SGmALbzJTcrvSl+SRpTKj
YCkpNFy20NpYs8wsyhgY3jx3gZ6qFmB76ldDtF5HfvH3Fr0ACoBxRI4ch/YMqDM0
17DKLxWb/jAppZC1VwIYeWS+0Wmb8g2g6h1ACCZ0RLD9IADnw9wNt6t19c7Lfupn
VJN8F+aQK3NNM5zJE2mG5eXCVEoxAT/8ZvFjALZb41pyi1+Pd3g8xcmjKbdejjGi
n6yLGdRgSgA+yurqrtkPnalhxSCIcAOCDdZpAh/Y6wOzyTQIKtuOOVrl6MtM27eV
kBJVU607eY8VfwEAW0HCpMa+lVMqalY8NpQ0P3C3qHDDL/bu2wbonP6wrwcLFM95
CMf2jkMD1jklA4IBhy4XvIW+2zfiWVJl84/7MQOJnxbEY5duzdCSW/KGreBbF1fX
pRitM++W3+RO46MpChlzLFhpx/kwrkv9CwDY4+w+SmTTqeQzkjk85iBoC+/Peyfz
HxY5Tf3tg+FZMRWSPzqkog+YNUrKwx60BRVM2ydj+0mT2yhGGvW7vrD5w5VLoQS2
JJ9px7e3PSnabWM57urnZYRZFxrAAwf086bUn7zyXD02aVLKhPoxujgDXNvyEIoc
0MoQqmfjYMTKMMMWv7yMURDKM2+jv7MPh45qllBAPx75jo85VEApECVjCRZDXcOY
FwwKEedTEqf242bXOk2nwMvBnIMiR804hhRGh4k97v9X2WpWCtNASUbYIWn0kdvM
o175T+Oe8cddUpf9k8COHlVavNI6koceTYOifo+QQBupr/0SlEnJ8NKz3hKyXvu2
4g2mlNPLLqmwnC4Ru9PoB9Tgw9vq7dhSh5bQWJgi44q2j6D4Xfi/AC/GcozuabJj
+KnQHRcRtBVSbns0OTkAVh076nLWIBUcpZCpB1EQqKIpS4ycXJOeYLEUUFtkXqUj
WjFXlb0fcBM2utu79LzHl3XYTMZL4cmEKazQdxsqqJYUHWySJ0U8M+fwKO3lKltf
3sKqt2LzmnGl+KGwgFBqgxxJVp9n5CdaKCDM51SC/yMr2vmD4hzotBr8LZZd6Zl9
sj3s9LBN7dRUMu3OdGrkE1NyQKxd8XkZgMo0+DNb+5ZrIsSmOhKYAl9hLDcl3O/Z
ncMWHfSsomFVfj4h1QZ/fG6LAHfLNmGOOwDHbmb7/DYaQlQG/dVCih/cn2LCRO3X
zNsoBgQzryJjJsXyzKsZ6RLnRugOXWjqIE0cO++JnO40RJ2Cr6myH9p7e6SJP94R
E+TtKfynzyB/u7zZ61woZkG580iMUetb7A34iQL9C2iLfjeePkVF07YQZFmmyYI6
dbFjS2/XXt+2oFRM3uhRQe17KOBztE+y8WEuxCReFOiZoMsoakJl9s7jZvsUdF1I
wz5fyXKc3Hc41poVYI6tvxGuQtaMN1ZhDt0G1glQQ/VTYT07jrY3b2hXYoLCU4sK
ZqRjGPb0ec0k23SR1qTGhLs9LFCUEjq0j6BO+ZCCQCDUKS3+wtdeW/B/ir+NmCz8
wWcjGbFVVnqa8gV15aRAbOZQEvHLEcIlqB/rG560r8mndqo4zVRfsYm24dv03ZkQ
q4LVBISfb3/2EQVBaddS3O6IvxeRv6eoGf2fNF2Cqj5Q8UbmihwPvzYSMyRf6c1I
4ucEiP80A8nzS9xzk0jGGS8+PBVUnLYfcdaNRvYhgVnHRzDBuc0H3MAToZ5LRVh8
QB+wmbSaM87WwP9y4MdYQmdSRR1cvuSGFIA0Vtl6NEiVw2nnFjf45WyJqd+TAr0n
OF0J2j5YgX8DmZ5TsWJn8XUBER1yvOJETkbu3m/eFakwQPWLRg+cBVd46By3Q6lE
hg00j3iCkU6R5VnXw5GXodmX2oXBEmMbQv9RGJ6qMu8dptjTjxd8/bwXx4SkvvJG
8NfYnM4bmIs0ZF1nASxuzKyenxtdfT7RiyffPE7z3ziJ7ouR7YnIoKiJXE0QQWFg
b9zx2jKnpvatmgyJqR5CP32Rb7kltEMfKcKoTpa9L+ZvPftO9XdPDgkhnFlcvg0l
q8GC6u+uAejFnT9AxToVVP7BzIpfkEVPqxsqzNWFunV1LaKz7ZU21usr4LsCZVHJ
y6V3H9idhx/0YMkeHy5dRWirt3tqCthkW6WhtcRYdBCciNJ9hWU2VUHLaz0PAS/r
BCi6Raf841iXEkJ04eOU22NWnEGaLRmsljyHbzjLn52gWOwVcHfxqRhBWXpCdGeT
ExPSbykDy5DV/WaEfAnpIulbtnLuOp+URVq9OQGGw929e4A2NsAZg1ygqfhXEqec
rpBxVqthbgS8FDEAnGlJdz5fLiPaI6zp6Df57W/eFfQdc6LK7dvBJCMAQyyLNVi0
4anBkCfOev/imR9HI7q2qz52DoZRqQkj5DGKgN1WDqZeMIvDN9Xl0B7gskfE/AxX
ttDu078tgu59kPLuXv9FmTeuhRFBvhfsn4v792jDFfaoRA1gFQD1Yj5cXPPfcHKh
dy68iHMGi87oVCgL4wgmrc+S2VEnQre95NQ3eoWAeNktAJ1+w4TlXTps6cXtMy6g
h6dV5HaU8xlfux6LJAX0bn7/kmqJAi6tRkqdhqV+Qk6+Xx31/Vwub84zKynTdwEX
MUhA9adO0mb8xWvR7E2dtEuzGBZrUM7scMZWvuVlLuDGMrJAwuqey4trOgG9WlpU
ZP10XessoKt9ARfLbGb5xcNTfgn/M8vBosbQ6+R0H3J3U5kM4YgeBDoMtXsPeDig
GFIcf0YZuqUDJkwAAVVXv/D6kC3pmiV0FLYFzAJUKg27FKSnbtWv0nFRlC5bwjV3
B5JMkVp36I1mBOdlk9mCTXmU8e+49c+Zoxt5oXsVgkpSs6S8woS8i2wWZ9fr6SVJ
xclvV8LSuYbidUlxyE902qCAdDGwa95GuyxPH+CMrbQooopM004lfHDI/uUPHygs
OWasJOAVdKPWboBX1G/idULhkQB2G9GI7IVW+ZqsZe/ON27EB3/MYC1JPV0Pvgp/
/AWlYaX8c7/8xJOh6ppy/TTQIf7U/AfTcc3qa4CZBYmMQKWJRUumXsMf49Ua+l6T
sbF3+gzJP32xf0xCRsv5CXelEqh1XMmDgYvV5vrN95jvquSsw3f1O4kjYemh06PM
pCuS6VHwOU5QHApWz4C/zYDD5Z3ggvJtykyG0nmB/oXjjSOlMfebLYPvkhI1OFO4
5qXsQDhL32HDNWgyRjyrHkiLmQJC+dLz1G9LytM8GsRWj+fR54gbO5cL8yAUWxCK
mZuv4mEySK1SBmZD8ycRoGXh6kqJDL1bnJ6K0rfj1idQCbXaJjxbbaJFE+bAwAXn
IK/6ktWBAlYdOGoyTikxwCOQnd/mUTLhUdsaQXkEfUVJQaIdZ8Cd4OnD9mTXV4SH
OyfoIOejPfU91R21Zk1Xxsit1SQccipwlW6w3vo/IxlRBKdDd0zekjF2xHa8dB3a
IIWRsYTAHvHkFKgeo18nyacKhyUpCp7Zv6dNWEyeTmlsKcfn+D6VxMAN/W7boNPT
kcd2Tfj7dHft1UOJ6g+vl78NXett4frPOS7M4uHf/oNu0ejrqSdt7uB3tccVR00V
LOw1sICK4IhUpwJB7uQ5FkXd3x2DO2fS2k7AEYP26xIXzFuCAoq1DjJCFwXf/Me2
UVEa4ofyRAFELpE8dbWrh7026RgUDYLbFWKrCKY5pjFBlln8RRut4xBbiAmBgoRu
OBFP59mCm92VQYf/b2+Wtngjl2u5ZDZDfJmHdWptLFQ69BQwQU7EvtwYI1x89wlP
Kv5ZUig8nkTVX4BCds+bTh6NtSHHuC/psEyAa5DE6aOMgAXVDszs5uKB3aSlcz2W
qpkky+nmo9ky5apWAq1LS4tD/hH+N6n5oOoptYJ0I4WSoG/EBofiq61f5DVkVX4F
uLsWiB0vbRnvICpSI2KI48l7kINk7satUs09s3XlhyCQhPPe+gZh29pBP2Ckiyc7
lKY5BPtpLXJYr26p8l73NXg+zwEr4kgAEjtT06XuNks7Dv81zPIeng0zJvXBaqwi
0nSADGPC1ikf/0QwuH3vTbLCA2zHOez6ZE7VIBH7G3mTQE9Th6XISRMzxCCf4rBy
/ldgQl8XkMGLxz4ZXaNf+7waZ2qbfZo4Y4r8eDDtBlnEXX7ozLOt2hccOggKOxcM
FjUjFCPePopOGvN+Pwz8DX2BP1mF5mdQAIolrvThWRPYrT9YEZAuVEOFM4HiPJ6x
WZsBfOK0sZ9Jfr+c8GCxZpwDBUU6jZTguxWjmSyi7UuFUIlYSVgHoxliyZ8qDbtW
hcijkIzCzbFrccXxCb0aqRcyiWpE8yE3W3RTZJucbJzj/kSsFhuNl0Vd/GJlEvmj
mudLnJxb9y6PMxAGJ6gtE01FYZqh9+Mh8rCOHuEZMkZQ5HJauR2zZYfEYuwjFnIw
nUKAKVCivNwsYSFITl4dXh2zXASbs/5ABz+6Tnd44a0HYGlDV8HBBLgCUpwCC0wK
EV6rOm3LWqI2KktgrbdMoAl9OwhCBX90+EmHWqTTC8amTtPruC7Ruy39D9uel9IL
C03//Qqyx+I7lxs1F+g+iB+hWSlvysKSJ1RgNgS8JYxld4o0yl6YCCs7UdiPRvg0
xTva8MYCcjw08iMyuuJVXSC1IrMU83fAFGQghuyrTBFNgpq+TCV0E3a9uJ6Atna8
uKeLLKfR6Ko2zUkuhHx7mo5+ohgKqyInuTR38tPOa+8qb7I4FUFfMyPokfrov5Nk
wmss17vCO7xxD5kZD7VUjGjg9xCDbtsrlKjoCbt99qqIp45L0uFE9+wLTvHe1pgU
B06yaOZB939FePFa8IQXSTY6hj6FxG5IZ9ry2VreQ23rJyWiLOGg0VxB+LYokEB8
WuY8qBYZJCZTFemv4qnCQ/R9oEr+yLRvm7lcP0PFKeb73GJCF4WjECWwNE4EBo2i
I6cT8evxzzKk3+q7k6K2YQ0g1EBSE2huwY3SQEv3UEDz/XhZdjm8r0oB5Htre3F5
5RyI21roq7iyWI8qdN2n+kDfrdTH0OHLj/OBNk/7DCtw8KZj/DVNWN/BpqeUQDSU
M2gZW9A3Kp7mB8Funew9E670j8I8wVGDSbpIub6T2D/XW8A/zlqdFJ4ekboxFeZR
p03r250h4QrLCf1sOY9Yk7Cu98vF2Ow82fYfWBCikIVdjttwmk/LGiXURt7J8B33
RP4cSUVLTsWtu94zTjAadh1wyJpuOa7FQmQKQoYgEFgJirkfzQVhDBKoeEZyQcns
r1L/1b34pkurETQ+Tn53VFw0K0ym95WGxb1IF3/vgFln+Byx4tvZYCj9/5dVqxLG
YzZIinvc8INdNvbwFAv1oIqOQ3RjcuPuen2nI92VxCoplRZD/BFV123+deTRHqOl
dP/MmXxctacJzB+MNxh1+ErSgeiVwfydKv5OS1v5a3OU1zUCk3bbhoGoUSwRiTE8
vhJUZ4kGfrxheroTOfAg9HjR5yywHbSSSklghSBx+2Jk4EI9MZAfvdR18dDXMdvb
3nqlrFwelu/vEH9X3uSpit0xkW82Z8XA4EItkUZup19gR0G6MG5kJfFLhCZ/Sodi
RBbWB8KROUT+pljWn8b4R4OmnZwVXyzlVykwfxPfT721KPkGitCgRP5JevTUSviJ
XIxNkZR8XOMBDFNZhXarmSLqdHqUMvLuGaMWQCMsMaP4vM5OUdqbe60IzeJLfmKX
CS2WvmjN+8Kue1hrUdSka9kCI5UNTyWV0JosLq0+m8GJtecB4JXj/uW6bReAFRG2
9Bri/ldvEG69xEDFBN08XwP+a2cvS3X7bPmsVT0U1O7zpaQ1Fekc6f6k8SFBqRBN
JiUpuAfr0piNWMIdQboSQZWGtmGirej0c3et/i1Fh2qq25B+O0iM1o9IoEpcX7GL
wpa+IpFwMZh9kLbDw+kpYtEPhhkqeBfxSOrWbLVG1RgHiMkhcPSosXZpO7avD1y2
uQ6MOrfVUvXviVaqNbDesSC56LBVZoe/qA2MIFK8NS+hsyG38f3oKCCmVz242Y0z
FQxBtKj/+coI7vZ84tNkrqQ53+mYG7n4vIiUavdT3C1NHTD8FiRow1H+OXoP7hZm
OOD8Q99GKZqbL8obDNQHT/Lp1H7CNutgyDB9wIL3a6DHL+oGOqFDdrkgXsrH4Om/
9PmCgAuXRewnKNK23kwqnhOiryJMgTAnQs12P1wnZNtG2IqqlgjYTsKX2T/C7/1b
I3tWltkMEEO/a5DccIEv/6omp92jb2nm6U2umjsIIKldJr90KVJgEz/bU96wQy+V
+XYzM5/56IXinV2UhbvabpICp54WOY7n1Xepb2c7yzN9ueKESZCrlyPi7/bugEyt
yzKFUOnrsgsU5XF2bRacB/j8vM0hsCFaxQhvJmxYkgJXDXE9NXQOYztGbfy8tfxP
oW3XbUMo+EyShthozTSPSaawDIhDbA6tMDNMwmYZu5BrXz0DOPW2Wy6lzug7Cs+D
xAuXB3pWAP7NsfUP2vBPd3draHieC+oM9wdC903zFhn2d4u1nTC/lTNtpXhsOTGT
OdNsPVVOKz4APFqLbZlkPYIFVsrdlADu/DP8e/1WQC4pO0KP3ApZONARO3bYzH7c
BaM2MY/4gAVo3H84kHpME4w5BYPZoaLT/iSbgkZ1Ss07LHWKa6Kk40ZOR52Vec0Z
+oB4dX+e9AElKs0mZBJe84TbCGqvyteWrPNj7/kGa4eLD01usyBCZVStRI4YdEmb
tsxoK5bixC8/shKkpkZv2EYBTG5zqXmxtsMA+ELc2qGIc/qUx5nvzh/Yz3hHfVk4
0ecuCmZLPvr4LiXtZ/vFYCUE5Gg+9tgmW693NjixaJw8W9CW3mcnB0DAZOoEKJ41
18Nq08643v9xKROdmATzFaKMr4i2Mtu03wmAj6uvZPbKa6Lu+ier1ckm/FVvlwqZ
Vl9OXXDPce+EgbWBkiOBIxNHRVNU0v1Ia8QNaf3KtDn9ufe9he04WPEmYcc+fAE6
p5IFoHQNBBXXZeRk964GmcP+xFXk2WVhI98Xhn6pjV+pPia30FTB7TXiKRayZmzy
Lj7X0R3t81cqO/11/VLPlt8XGFpeezE5lMTYIFZBK09sH1aw/2QSfztXgBdReC9E
qFDoofUDiIqNKhtVBt6IUrXaSGEd1YYtJTmZ4Ocjcb7ls3LvYgMMIZlBAGZ4p5vx
EWpdOeyQdr9nfWt2q+fO6AHF++VMGzBILWXWVotz/GPoW2trmSm5wWOBuKNLGJvc
0hsG0g9j2/XSh5w4fJIeQYO9QeM0jguGYpDRkGM2PkR5O5vKTvGYUYHZabtI3pqH
bb2AwzZ6WhKThy82E3IFWLRKOug4Z/Zs85JHVslLfyJv0cBdH3i9c3i30Z1IGL/O
jyi7TBYNc+IIBpPGZOsvijpUq8cZuoUFgtLeNZLNzFM9gD4WqEoJVu6bf6Y6l0u3
3rFh0QTw0NM/5VaI/6GA35lFVqKPWVN2c+MgIZV9EQAkHxQulHbKp4xZfY5dIS4f
mvnwhy7UEAEIueMyRg4+guoeK/C5x0BZLoG6N9YndqQ2ZSxWm+PI5um5ezy2na9d
lsuYut+UD/Oq/u3DXg/x5BxghLTB2bpLjC0FbVYmgZYCbFDKlSR4S8xMNQm3QrKa
A7FpCBZq9G8beiIrJNIyULNRxUlUTffSFtbJAYqr60I65T4sLP9WH5llKlU4o4rC
0BnkbgqCvjXciM1AnYyD3vlzozVgE8ssHoyh83qsp4oiRb3wcawz758Ih1JfS1MU
a2JLjhF9nHoCLdmGK398GVqH1pIJbUPoMalBwPo0PejTHBmDFkUrmOKlR9tz+a8h
l6xHYVEO08NcPgPNmaUreQyglx9rXzmpd2N+NyWn4GeFf3ZWzGdFTo6FTMXICccl
3++QYMNGt/Htuet/zrRVLRqOnaUzKoOhgdn3/aWITXaC2ZkG1/rODgNixOu6UC9b
QDBTf8d1KzhuTXOhTduD0uMwOz7a8UFFF7qYIArvfK3kJQuCPvTQDxMCxNqa6nkA
iRewTM818kQYfooNUjYsnG7wGR4eV/Wf8JcD7lKwGpA24RhMim3vKd0LWaWb2RNt
YBztJCB0YsQVQix+Tf9IKHuKWfsG7eGeWlczBdo3EAD9fzeZtlmwwYLVCdfB4pUb
hYs0DLOWg4p30iskeYBrkHz+e+OJ7Nyx0gJSViGOzqTLHYeMV1ZALKw9SlhKVvan
4NI0N5yVgjpert8zAO/EpNGXAbiuZJptjWQGdPN6n2eiSA0PADPYA2GbhZe+X/xx
V3svbvKGBmo9BbN/1m9JbJCDhhIenyJtRH+RmGOm/R4XZOg7TkjUIix5UYBrfQ1C
lWs6CxKDoJ1f2QRuMiXKSO52e2acKV2scvs1TxaOJ4i8zFx5loMghtVwmrfK3zAS
Yxsw6jPk7FSOgFeW6pXeEWocgtpxRha9JgLEHrDo+EuLPYGPcYMqHuW7eWGuGkAV
FCP4dYWXAbJY7zCa4x9cvp4Z7Djd1OC7Z32OYxiR3KPKdgDCKwIDajdbd3Nw5ny5
jH5Uh/D5aJuznvDCoLE6/i3hI3pjD+RaZix+YDW7DJ8gD2mFYVniKqn7/e/1+ph1
/ygM2tLFUPXtzTIJIhxQvRB/ST0T1NS6fTH5+MruRr3PaDt45H7SO77Csm8Bwk9F
mFNfkoDWZ9+7R1yLq/PBE56VVq+RidOA6liixN/3QZpjYphK0HecKt0XAmm6jcYb
oGisklO2CY8RfyKZp6X5e53ltAtT2d91w5zPxlRm8UteRWRb1CIRCqfM70sj0OdJ
fDw+Pn9tMHYXdcKTA3zvLIGRV8pmzxKtIVDujro1zvq6peeR31xnwqFBT3WxJrDx
/WZ69VEPInzfOcjAYJqzJ+MXEqEIWwFkzg2VaTM95ZGRFUi5sFMud+oJUQbuUs3S
MGIA+3jou7t0K7mWY2XSLnH+86wCCXLErAJxUZOe0sRtCJ1jKH+KAieUplArSuri
MsivyKVRDDpN/sUbMKpupSFiFjSPZOQRgS1a5AJDbgEfUjdm/heH1k6mqvclMp5R
NbGozRX1UmXJe4lCXqFDgBZO1+PX0UiqlaPCnstYRHH8j6U74dT1eMbx2kHRCwVE
Y7DffJ0FCkB7tjhZ9A3SufsrOtos29DW+kqQoXrwiKg4NaEafIB7H65Kr6qkoBD8
WxUUGCO1OreTepHUQHQFWrbh+3E/bdpkuTc9xkITLATeevAj6NmdJyNMb2Gji+HD
CcSg3E8ivwXdwFytx/03HGLE30jndOXuO1UVMm4yUUI5IKt73q9iTqJRmZ5/qW+r
+9Gf6tXS4Cw6LHnEBXr1lSod5zXoKlnM62vUwvR5XgyHF5hpK09Mbc8W+UogE7f2
GBwTLBjKtKzLnStJA051GIgR4yC3fyqsb7lFBcrwapXe4wKDf0gM38+JRdngNS4w
zkEdNdYGwDKVTfiQX3wHsv28eXY6wx5hxljIV18pFxEW3XWy4IE4g+VWNhOkGBMD
ArxbYLCwCWazwZ2Tj+yfoiHFUC/PsG0ZhNCNi5mSdz/RKyEkPUv6X8DI04XlRV56
eI138YbOCR81ZgC0EXDWftVmxOVtgVEjcyLUw1FNv3YmAvwDSXjTH12Kz6nu6qdg
eoLux0fDS0IefFXFXMYdzF+VPuf20APLgvYnPIXWii30Zc/Bk4FBmy7nWadbXCWC
8CXkyeHNnmzCVjax7ziuMP7MICjPf1xXwYzp4bbOj5D8uLcOJcD3dS9OX2f6hTbR
v5qtmOOA816Y4qyJiHT2ZnXVQlTfgRnBMalIIeLNjTMXpiIU7B36gpgjPHgiQrih
uyww2cM8CIKatf2S3s2f7PjgCmEPUecbsesYQJPKIqTTC7KTlH22sCOSTT08Un1q
Uo03raUoWiVkho/E62ril8wK10JxvXVCHmpDKNr6QeNx4QwTMtzHr1MsfvP/dcvM
eIdseYkhKNTSAkU6IBj9E5ZB/sxzKUgYcYWIoH+aRG6FMenAexKuKQjLkyt20U1J
bFK2qHuYbM7VZYl/NGG68n1BnaAqL3hfok19iqa+9mRuN3dJ+Z9dKi/ECN5PolSw
WpsSyyl1S1OLeh6x+KDC4WF26zMxeGJqStfCimcpywt4XHKYmmeBLYEWyfWJsqaS
Y6tyZ9DjORzj+O/xKMakhlDkT1QmWkRmvifcObRbs8IfNZrU8X5ECsXMoaMVr4Bj
YQHmfif5tgL3DFl5MX3Ug6VYiide99+X09C/H6CeU3SuMmjiB3mA+Mbn4pon28B8
qrRv2Ybiuti65R0J+0LvhqmTXVM+z849Y3sFm4DOu5rk2t6VnHxTX/quYV2xdhfO
v8us1XawByoMMPld6PCmaSry4s6PUa51R9C/mfiOuMrqmBlL7M9sDRyXQjKBIe8H
fYp7ZLtxsfjdI9jphhC5IpH87Ow+Mbrq3kTgQpMwEV88beGZawFllrLqxF0ajQqw
mQy0FZRbI2KkPAXWAzio7UEmFrPp9iQDrwQOfiwmwWT/Hl0Uo2v21dITO+9c+BFN
iA2CjF+pomGsjIJI5+yUhgINiO0LcO8aFrRDBdP41/XYvgi086JBoTu3h8oPqz5J
nHdrgKBr0SErg5+11HxbGiiiVjB+qaOn0OcSQwjTDDbc6FiU29Rar4sbm04sN6jP
dTvhNEvxPxXfKMWd/wXti2bctszsBI+c9dUj1MGINvrhrrv3jlI6a2xDaSVvdX5F
f5rADLOsLVRYK39hodoJMTsas/bP4qlB+K/gjSLlLrmtO8xF+w9kQ0u/iwNnWEue
k0NVp1KO9uWFf1gm5KNG2NCki+Ij4kptHvwR+qcXdPfzbChNwSQKOx+nkejApEtp
AYehyA2jHE1rrEiFK9kkauKonPsIZSPgKtc0HqRYCaKuEBrjwizexUOoRbm2knVP
FrxJmXlfBOFfpGf5HBt8hdRYyaPxZ1YbJRjiVMhqnxVTVT9MUwSxzTyJdG7tWGsf
jMFU00tH0mNFIeFisrarPCz8LQ4Ur1PCwHtT3/1W/qiPi3CtXupjOZBUZ6xkvIdG
FnLQY58WwneR6tNVQV6qmf9j7J32AFmWKqlhcuXlDAeh73Of22Cmyeif0yI7C0RU
+u9Vp8E+Ip96h/15ie6thXreA2cKoXd2pOxf7ZOZMHAAObrw6JNeP+W3WmbpvQt1
Tl3UPO6UT3+6609tDFKWoq0PDI/C5E27eEleubq9hZI9PXkJgH9CCbdpKlQTZzZ6
ha+VowLwazKrC7l8Yytji4VGDxx5S7KYiPTj1qoCl3ZxeAZE5sylTcxNWRk+1w+W
u/55G+8d7SV2hMnWSmQRM4v5PJb5zZBlcOR1RsXuulD5TviuH8RZvbwC1VxZV/IH
COjUwsIZu9blccEZz11ddoT4yZDQwe1Z5BxRF3MJWXmTdwk0eG8xQ9WwPDQHQsb7
rRSouW/RQeOgTVyxhoJ+WX9QG2coNKWZKatXPjf1actGvYLlXN9kQG4lALWNgSfE
1uzESUocvUFKFnBCBVUSVSeNbgcIBbD6VaF6X6fBfmOvXKMRN/6VTCVg9iqJM2Na
ovl7XwfvP/2SKKuAan4qJSLSh6Uv6DQTHkVbkiMAaYCNlnlzQXmAqIbe1F9WH9I0
vB1ymAJSUYOYt0lF1vYNNIsIK+MIuXIHNTkZ4aDEp84Gm3+k625LKRBMgnYuR4MI
ofCYD3xZdKD/Ks7pDExjMHOmBB8IJkxpZz1aCqmfVfhhgEti5EaDOlYxTDOGZZ+E
6B4LypwJsdKgzTWCGeC9RWYsgxxlnK9X9QVB2oLFDBeVWl3omqRk/NWP0zD+rH9Q
zP+QA6tB7bbJGDW+bPzyo+OgJy63n+tHE/6diEgEFNMqoLzAlVrseQptVj4CnED8
+b4v+UG3vmxJD+xvtJSPLxvQ13+8vvz6wRkmaODaZxdpBo4u7DC67bF5dzJa2iRa
YBR+ySEG1TKv8OwW18UtLRMX8g3JCZigsBCzL1z+esZJ8ufLTfHiZ4zdeTUkilkl
CTZ45U7w0ipHTRTJGqG3sMMnWtkHOYQyAHlEqJzG0QhrOTdfxtu1l2GJp7MlM2fD
9l9+oRV2KoikgIUhVCNo94QaiAMwCBEeTn/69ImfQndlqAQ1utZREIWJ2ngM01CJ
2CGEcEXIURf6+2Ebf76QMgrmeIKen4JHBaZw/jkD9Yg0IpODEuywSuYf6s7Zf4zN
swXIzC8KahvRi2RGEDW9Osc2dYNtJOFG2IL7olgUcJ2RbT9+D8F3jYnyNzzzM+Q6
ozO2unpdLWHZ6WqobN9b6Sed0Oc96OruG9k+NsMk/RWGOrIWPXiEnUhqTN7JAa8K
q06Nf+mtHnp6WykMSdPfy+QZRvAgPfEWZLovF1bJBpeCQdx7ZEmTmTIBVnamf76B
xb28WlkXzxlX1LZWyUKzPNGYMlkA+CQt7I6bZYO2XLYQ7SR3xFB/RTSRwceYEHzU
vXoa1QCK61mVyCQfqEOd7kpDd8PqtS8UtFvn8b0Ac5TRlmsOjVjR4/XRbqCOnrbD
NyGAl5QIQ2Yo+7dCaEK6BTh+oC9BBZV01uY9L3f+LVbQnh3xEGg9W86zh6R1H09v
lcO4nQdJO4PjpY1dLbUlODbI9DwWeSgsnWFRZriwswPGnHUehVttFuvnBMbBTuzh
mGHqNDqiBiGXAQBdkPTg4zG3hTiVM7+fvvznDQ3RtrtWnAvpl170j8rlIqfdCplo
CVJBpcHeIf36GFUOik2Q2PKWi+01wmUnv2ENlD7loStTB/itn8SGVLjvwp1QdHj7
W4gRMpiBklcX0mJcFZjOm/W0gExvT3lugDwkjyGks6dMFvQNaws/CfkE6mWokevV
nB8g6AtRMiu3smEf36nhLAsOM/6R3+qBWuqPTu1TuGfJYLmAshXGBFPvVI17/XhB
WPUm0NK4S9UmWG1XL5hgYtHYeGLCUBE+qdrcSrmE/gv/hTOrFUqArG2PJ6/7+qDj
zYitRQdPmOKbigIHkSn+qMZfX4Esd1v/Rrsa2Pm9LZ3KUQuNbqWnijMI5spxgkFj
heiVDnih2Hv3BMreTsHtZwAB+mBCuWMC+DSbEykiLVATCpKJGnFuo2VQpl1Lja6G
P9pcG38BzBtjojJ2fRCykVYKzQ1G+BIl3dOU9ZmSs/aDaBLXuRfRiLcJCT8prUbe
Jj9ZESx6xZbvC01W5jyVmmOHRbFDXa29h7wtpWijaoscQW5Lr07sruLbTIpmGv6Y
1P7KePabmLUFtChiTTia971TsZLFdj4OWxGQ/PHXb4gqRP1KB4miQQRJ1ENUmVj1
a50tNoyLR+dagbNsRpmJbQFLmdDfzM/F3QPh2v5L+K5Tyi9H9+0qM6Tqz7iSm8n1
slTh+XwkI4VVVWzEnN8TrZip2are3AyEnq9P4T3duWEx3rIrUmJiBIfT/ZjX91yg
OefBxoOz830eBLCuLbyvS2+eW9N379RVf4UPNPwA++oCbtUVjMSL26Gs1HiLebNL
2RGtjL/MnFRVHCXDSNi8miu0B2vPemxl/W93PIstF0bCYHLM874/Y+XiysYg9Kpu
FzRBO7Z0391HJQxKDubJMQtrA1fdaP+1zp+6/w1WNEFg6TFkKOadgRCVZ13s7dod
3Xd0QRVHFb96nuouSk6ej+bE9oVf6HelUPH5yKzDX7ArvE34NaWPHay6lpGB9clw
d+f8hsTaFOTHqC7jaB2fRVOLS8XXV9T1UD3qyGY1DTJqPQKJofR9rEo1Z0+hyTiO
3mrapwlXftilOyQXxWl8qUZ3c/snE8iVYxgSwPdgUyUJNsJP+VLd48xtwycbo0zP
SCuvmxoQ3lgaJG+krrvGUmxn13i9p34H8b1SJsD6pKln3szYk/EXBKGCiwqLuWdo
y9rsKz4Rw1pi6NjmObaLBynhGO+xWeolFrN5y+g8cZpVHqSf0gLJ5+wt1zU55vHe
qqPSQSUGCtAbAT5ZRQVjbXoeKW/zpNgTT+gWPH3WwcuIZRtMYr8kJcUsfHCO5NNw
dDjfM8d1+3dgnO8lxd/QaynWd/ArJi0wJ9PCXNWioOjS/LtAoWlu16t5K1JDS9Gx
r9QX+CH0q79yOIFCRg76yYt/IQmTY8hp5LmpCdJmYX++KMTg8fFDUTq09iFQiQ1h
cLJXsV7MRQ8SMCd5yzhE1sYqabXHhdwTqCQvkKwMcrGNz3KdICanqH3Pfj3LLIw6
ceELY0pP84NnoSCiL3JLbVs48RaU97c6dVyNmiRqIKNEHQgzwmHfGOyeOLZK4Aaf
/ltWKFCYKLBI0LhQP9sTAriI2wA7an48TCojdYOrosDQkOKMzoASaenLTgbXpUid
s7EcDCXGYQMlF2FG3MwewPHUYSTFd/idxH8ST6QxbyJTaeJkRPhta05Pq4Npvz37
jMOw4XMDcM3084SEM2FJp4o0PbJ5xHcRODbhWXgztizZAtH2g0hp+I8HwRECR56r
czVG3/IFiP98Vk5ckNxmQ1e+cfPK/WJpCSuOZIlWCnuYPzxpyMdQuPA/TQWOAFeQ
E+Nv2SQCgFyEFOv33KZYDXEMMQpc3H0Av3x4hbu1sdwoa/gJ80lr6/QYiW4Yt0ql
PQXcOuWoiYhD80syJrlOOLyDDxmnQ8hTyqTe9mOelg6zmKCwxgyXYn18mHv9QlXq
+M/VS75nyfSRMju4OW7kYgdxcZPUIK+mmnWHjtABJcHowlNtppdcvRT0aZHHRwUm
rAHRYYYOdren7Ie9ZIo7lrkFOWz2dkK9ic7ffiGFozK3KUMOBo/a1c3kgaNkOAlB
//guJejjmtTcsKb9HVjW38cFJEa3qihiWZ3eEqpq5UbF8nkYiTX5rj3ySYcWIbLz
UVQNoNl9Im8MrfMyTn+c/KSOlWI1o9zcE3Cv3jW9a2Mlu2bWDuVB4aRzLOx72TQ+
i9L30zi8d8UAvxIbqZts2fPfEBxg0Q5RJ3/7br6/7BHsLVgVP/S2lQ/toXwud3Dd
TEQQMKubh6XokI2w0PCq4YIB1ZfrzRX906d/p1sNUDOROoLdcexvpVapS4WBPVm9
oVBx64jboJEQ3AcmW5yX60Ahg6KHMkqxpiwQVcYfOD+nAqtU0lxlOxnxO9A9kDKj
06Swcl/HstQknujnprLxpi26UVboRAD57blQYfIdwCqj3kqT4e0whmqOdKsA458M
MpcHJBbWID1P0JnoRXxJ0vX/POQKLjteQLMu2/rKB/Osa/fJmiHj4H+Le9M/wWU6
PC9IQLZKIU3iwo895ZhLGrjhCxsd2vo6YEn8EIh/2C52S5W8sJf+xWVpHLRz295a
iXrGExVviO6WFPJKG+vc96t2a9vBjYlXkc3cqXhaZSB68HT5ZPQDfc5G9UmWp0I9
EcuW4STfoyGiXlXsOU02aVzdFV8QZmuqLocE6dqM7vLbpOCvEiBj9uNittEnQRvZ
fGKTNwetjvdughsGuS/21HyPynj8seSs+xR94Bp3rywS6PucxbqhxVR4JN23Uxwr
N7fNXNZWMsVH42aMHoCt7V0sXS13dCGhWWxv6sSR9sLhEX/5wtadWCa6I1Yz+wqi
/CLzy1mQyP/CcVuywWFan9431pmb/5lyax93wvs/MpQe55w87cWVmNs3lgA35uPF
VkamQyJ/9zZEbHx16lxTS1DXEz9XCEl0E5sxtx1OJ6MXGpF74rqsUIY4lPz5p70l
RKcCQO+rFiOEFEPaYnRNjbe2k2JU4U5nlyXtZuzrQm6Seo38jqFV0CGz5g4a1/ct
e1tQUI0f5QSnwwnuPwdiEBrjEEFkV6dGM+FMaCXsf6NfKQ/QDUMMegwQ1GKgnHtg
EDe5wt4xFg5pzdJLYaQhYmSdhzUq97oafiTd3GMLWFSBOSBR2ElVLVXwhSQWxvyw
kCYiwNWtuzBY6ZCZS/WdUcWd2d+UHbZsskGGRi/61mxdbMYHN4IiGqvgijWiJNqa
xoM1qbwqO1NrKT/tyrZQ9nlHg1HUtD1koTYpM0+f3FvjGYtZy3UOse/1riUkd4Z2
EHRb1HZWxn7VUJvoeZ7HswUfmpAvIYR/evSgWfIUQwoAiBhjNgVDBzMaAHTrYcOf
B+jflrgy4h1etQcBNr4t8l9Xrkx73uHKgWIzRNVUEg03bTme9t0vQJE/2MbFs1AS
JjEcnhyUiRBC6MRKKPW/AmqkykqE7tIKs2vFBbmBtrrI7iDyqSkTjsjUNNZcHhH+
vi/rNxRs/vIyYHIkX2onNiTl1yhPa9wZLitfNyCpOaf+nvEyhiKjnPXNTt51u0v2
RPqug6miQc5u91KrdsXwTSFGT9Ibs+p8U/q1KH6owI5f05UElK5pAtkt511iaroe
YPU8geNtAfYOrhnGALQZKSYAFrO0VoxZNmwhmcz+nb4hdZWv5gVxa86HyXqafk1w
sNyjzsswZDq3vrWemAUSksvEx1IiRlUBCSre4ngk5EgBes6DquNhOdH4EiDs06mo
5NKJAd5GyvWuNcvsdrwiQ3uMDD1UbM8AHXrN1xi5tIxML/7gOnxexUvvED0VbygT
CtcdYK55NbBhATI8gbzlgHzMdvnlZ+Bytx6nmzZ93WlW+A3h6PHZLqwNS00GTWVf
iKVVWwFFnUaYNZBtKs4RsbPtcpCk+rBsGw2TeqBrrkwb3qRt/Jw8h4S2TWnlib6g
pcUOjyGOq/KsFpaRT71et3XI+13Q84Rp1P99a2+OeiS3hsK61HBikqKh+rlEZxu/
sjHjaTE5xJy09AfpFyRMWdfNKn8skksDH9Z69NVWdcjv1fld7EePbFFkYYD/XzuR
c9Sk/QJF6Dh6fi70xTWGVyfO+pvf4YjbvQFGdK5/dwAvreggsWHaTd1YgqPjkPoB
fRl1Qvracfdg9hQWM5dU2eNZQv7ziKH0lFjWcrGgkeCA78kQJpe4X8xp0W89Iz/N
NHUTEZZ/NP0/E2uaNI8Uil7pzZt+d6A3xR04qpynoJvAhNJG1GdJd/24cxCw3HTK
6+plwiTOQwO3tIAN8fqsw8JIloIHCytAZyd6E/ndJ96siGjv+fpZomrOLxVRNRUN
U/TfxD47T4afkYruT3ypxQ+i0M6uTaZwUZuVKa7xJX3q4i7gUpYNjJtsui3AK2Md
dRu55sFL0HleKtLS1D2rhjVLx55u5MM/MGy43nRt9rAYlFfplqgz/NWnsLPj+/iM
17gQFBhtNHG6tln4mpSBiieyAIoXzqkJHJy1H3K9FAv/cT/Axjw0l9l9OWyC+x+E
PsZC3O9I59LPJ42/sLkJR2QUcdepfJgI3wLMLgcAkxzYZqS+w5NEGAu+grjdytus
tF37fQNFqjuyUvsXZbUqATLEKZO7C37xhe6T89CV3/GWbl2NKXoaP2tjDKIUW1Vu
3tIrbKGiIELmnEWr+2nBvaGa8p2o6hbNFd5QfvA/8eoZj6vM2RB/neW2mnRcJuQG
B2Cf3NZhi9wkPusm3mA3Q4Ly3jpNgaCXsmTyzY5ikJD2Qo4/X4bXSHx1VGefp0LC
nP0Cz277EVJ3azrtKa4o7cf0kfwGpReC+gPvs7Rj1ZeSfj7WxxiNba6P7YVpmDxS
uXCPEFkZJ6bEfEU1hkHWYlrZl5AYHZGGiKcsDbVEhb/7sHANnxvjt/m/noZ/u6Hy
eQnPhcWCizBvmBX+YTRESBnXtjCR22r5HxRBOR4/7t8Z1fMH59z0hB55PKMQ0bi+
DAXSZcU6ZEkXzYpg5tc6HVOrc6GyHr/bGTtjC0wopEU2lTt+IGMbJ2J3oMOjKG+o
qHI3RFGZHeFkUf7UIbzMuqWSYGf9MUZ/H2bTTIfjpiNmRfQj/eJkhLiSHqLEVHLm
aeNgQ5W79QkKmknhyoUcMB5uhGtBX1SPEdiUWemEz7lvCeOgoV9FCLm99tPnJ4FO
mdu5T16uzsBHEJkcej+PD2gEqs9uxi2L+o6t3IMw31l5Qvmr1EbyNyc0KaltLvlR
lYm+4dbnSBptqtD2WMZwYit+FDxyLlYxVDLLGAIXDIx2zJD4YEaeopVZIY4o/anX
43IALQ98FLrro1qpTt0Y5KYby/BvKbajNkR7yHJlJPW7MLp5dXrHRDN75QV/OWsT
qqGQlB19WHghjk0tFSYnEp9qYnN5EcIYj6IV6XiGGUutykEvu0u/cK8nHksGkpql
GKzyeJkpRoFoxhro0tJc/7DN8P/r+qW7zqvlW6QOO5BcTDKnTSxuz4vTOQN3zytf
GPHWMXQ9FFZVc0wsOMaooEllKgQtaRq9euWjOeUfDYxyMVqJG/qiy1FIK9yoo6/n
cplH2i0B6ZKkk6Q6TUZrFDUrQsNubBOCazMLpD6yR4DsRvxb7PPhI5ulcVUCWN8P
D8M89yi+QqNvyMEPHb+5uodHHZ/p9CY69qB6Wc6EJc1eckrmvHOtpZ6zuIVxRNpv
bHcm6R3NIrEm+O15pcmkpWuH7hB2LBfmZtJM11UbBT663TVRmB9K87oNB+GUb8hp
VKLNdRg3+xeqFUXe7mcK0rsAiLPz55qb/PL5QoYjIJs8MrIXa+dmq81EADBOkapZ
WXtMY7KcxVgONgbXW+EPLSXko5i8d1MwgPcltIPj1nWej5xk+hrCvuyjcV9JzNNg
3Ero1Hg7pBoD+BtexDjTa6cdvU7fvXawA1RUvuRu0styuUTMV1JG4FchCyzkuRbz
wyIO1piqwFv0erqV3l1doNxNp58m6tSbOW2Mht1BXQ0W7mj6BR/2o+4o1q9sB8A3
OkcsivPQxfQdfQ9yGincsNFIlt+wyb86jiZ8OfHr73/shy0Wu35A4rrlq8uYwGdF
tcnUrOwYN1nAVySYk3qfefhYxdgPvX9m2HJCeoCjNSD0gYuG4y2fkVeOQ693QpAi
lcFGzEdBqgdFA3FpO+PcZK/ZYxR4U3abLRJ1jAzoXzS5+HIkolBYKTDS7sInXewL
Gd0f5bRag2Ij5wlGEgEgRyxWAiwY11Q1AcGEnd5Jil5zUA+wUj/YsGnwf1MPYBwb
RJ11HwJe/pAGJjn8IqoKZQ0MO6mec+lS+8py7lygfbDuYSorUGhyvBdETzU8gFG7
N+Qdsvan3UevYZE+WJIbmIqbfP/IQQeattql+qXgxsnpC81atJ+q/jTgH8BlyjZq
Cayf4NP+IUDcq+C+7a4YMXKBXXjMY/LDMIvkyHFJhK7mmufYJEol83ghNxo/AxzP
TIjKPYPx9UfT0s3aYbnfhncTI+e+I6pmZZuQFtdzrEKAuGVJVM2kHXYR/upqcIqS
8WbtWGnjlNWrAcX4o2aCfnBDZHtaWk8MOX9sk2irmm00HKM3OY5VyaMzFdnurl3o
sfWUfZRmybRl9J3v7SLLr55mWOI+ZQidCCFE7Kpq4K00uBBcyPZqsuEabBIZ1TVc
TbU77V/LYcjKH66GmpIm/tYAkhrIMI7AcjyWzj3uSkr6jME7j06yoG+Njd93ReQ7
XGMHiLlv5QTyDZfsJyUQg8Vc0tiJAgHJwloVNmUpKUn39Ar3BHkgC2u/E8ICS475
Fm2+OuES5AGkE4PmqBNoXJi6f6SkaYV/SPwt/Ufj6NfLiwaFFuZD7plrg5ZDF1rt
NM3UI7FbJQaaRg0bMDrAg5P0P6W34fVbCX7dQY7IroZJku1dn8q9ZEvtcpRO0p+A
oHZvlLykwcEnk33vEk1aTTOSv2nXmF85LLK2n7jus+Ps8gVyYR+j89gwWee9alvp
qY3tpdVJWnWJa9IrZMJSYV/+G4aa6zYPziPV2WreCgWFQKB9w13PMcmq/r+mH+2F
YIp1CwoS1BQwgN0hrl9ChMmXETjgCCvhCpZW8rPdmuWILf/Q3tRJ5cEObwPEAZg9
qCeAyowXmqjFKMISV0eL9zZR9Ua1g7cjlW97kNVgu+UrBV+u1XfP1UWE1IhEuJa3
3Y8PWV6JVH+NDx/Qxe5WEAN7FZiCLXqPuTIJQKc4MkQ0VRaW3QMaFoCY5UBAt703
xQutBjdy97SL5zS70I2mnF4Uuf+xoLHTCUGRtYARTnHDeCOeGORoDchW/AQe00Of
+8d2zaBoGPfgmPr01weyOnUFLOPFEFKStvNyyrP6VL1aXWJkbDkl3gGxM+FuVjkk
6U9tF9amqAW1aN5WCZuEMHTC1KPhodk6Zr9xRcgrtgqxm2823224m8RI/3TS5Paj
PkVRjNlU4jNGqoyyhYhn7h0a9Yr4V7fYeeE4LQ2OUrOfOAHh5lHrph0NGVvarh+Q
JL6cK9EmQtbltrr6x8xA+6H+rMXYhSRSpyo+WbZnoIBujlZfgN8tGcNmoY4CHx5J
50FIuOsug2zGIgF9rWzTfBm27j2A0uRHmaclt9yIWJct1zkVF0SNCTQOZ6SHNR0V
y1yDqllrtBUcvaYynfrlkFk6DSYlGRfZuJjVOAVr8ZNCthSrsEk0NDKdV5I7wWjb
Bkgxa5c5ubs4YEFPBj2REN1CYN3eZ6zuBozBvoSKqQqVuY2BeUEIiXvOD0o5Y7FY
Yr9VhPOIdMEd4O5lnBJ7+zt0lyfIW4QIvv6MyxV1nW9nr2GtvLgcBtT763Y55QUr
3atwNubH1JG78bnKvl6gxG0aUOk3Asn9oOqilIexAfxDg57h9ZDrZZBeId3n8yE8
pdq9sOlJvvzDc7zP7ocI32uVbd4Y0PkltO/R0eKy+2sqI9hK++pnEc1MuuxntgWe
dsz71FXwOP0NgV09v2KHhdYpy7l699h+Wymprthlhx6Mhy5HD7Ms5Hh0JCYpj6Ml
XcE0X5haLEdJNc+5FFAXLzW+C+2tPOdbLOqctmF1mVdmOiV11f8Y5VhCCJPFWxvJ
/LFlql8ITPANgpYwBuwHO+ZaPjUG5j5MwAE2FXcFXfKAlOQVdZtAIV+n33P5+dCh
WK10yIoiTvNYUaPIw26nwFFixwoRZtZASBViu1ALrBuoTXfQTmV281FgPb49UUr2
ELQPzqZs83rQDFHrpebyEVBMFlrL39LOIs5lhDUm02Z1ntcuz9zdlJkwZYbuHZ0s
zkZ/KTdT+jX5xpQKfPYhsAXse5gKfa8TWFEOfAQlBFsC8420heCxYi/6u4QUeofZ
NtPTDc3aaZ2wepu9FQ3V1rW4U7HkFkQEEr1csfYclF7J17CDvmX42cvdAK1/J2Vg
t5jArz8ArqpszssdYUK2ADp4QgnOMkYahaY78HapatlX+B/lR5s7ieTAJKDW53Yj
C49nfmaucGYkFHlahuX0enerohxOrBi1eFOEoeevRkqmOyjjNL/mY6ZHimHmeMbM
9V9UZdykxNu31/EWLYNFGxa8+ygkKIMNIGf7QY8yDiCLTX+htAh+NuYgr4Ns4HaH
0uPYBLYDYK/yupdLdNwm7eupMQXZhIxQ42ZHKuTGifbAYtpcRSjzE6OzjVy2zFrB
nkJsU4Ri/p57VHqm9TkPwqqa3E4kp3pjh+ewFedTBSueQBqn/KFq/uXYS5pBIo7a
P5mprIiz4JYtKLkq14ru9v0IsfQIsCsiaxNMC22P1rA4uhFT5qBkt1bliPOTm387
iqwP8u/JvO3Nc8xW7dMNwNHAVTTn8a8nHuez5IM+AdxBIQxcSAxSIrTwwDJeszX+
UVqWYu58gJ8VI06nao+zsktI1D5POfmBaGX4WkeE7aoGy1ST5pRo+91F/fqbtvJw
opfnqKzKSq//h50WwPrTpbPedFQcpCNQRmR+bCAZ0E9ViaCPCklz497uAJmJunTK
rKC9qgeMoQqsZsbxBYM48EJse3VRZaIxnV9+isIo1guGRcgOhtuHBUddoah+V0uW
Juf+lDiaz/nI+lHfp+JjZzBmWtaaDsTjitiFzOR1JMZEZiqP+NJPrwBc1sqhrRiC
vk9zAAX4LCwttLC/JvT0BJv0cajHQuHDWNlw4/PsTrJN/y5dpoi1O73EFJp8O3Kv
dPbUixiV1cDCvVKaHqkjtFfMI4iPDpogPub0c6nkr3/DGxpzCW2T8XXTBJB3S7nS
OWnGwcij42ywo6jtdfw0umTAG4+DNAoopQKCPZKy41LyxXiKHaT3rTJbll3cprh7
kWtJ2eJkR/JyFU5rJzlX0ByFKDNuI3nRW8XTDz7w2rJiTcQEUMShtK+Xx95yhNTJ
EMOS4ZNDnBERwL5k31EK1jmUITJewVDSLX1rRvoaQd+VySZbNm0Z9jdI35jyyh0p
gZu2fHC9rDnz4BO8xlanVcefde2cJqJhb2iv5JSbmFv8VO5fwjMoV716LYL4k68z
hTwqwKv34loL33O3fSMuIK/QL2xt7TvTd0+DE9Djr6xx9/nTJhl0PtsvlcqeFP+z
WNDKoz2W6NyolO/raTuKzEiDdIwneTRbIYoy4kmrEvkEzG9zc8aC+0dDYEAuPI5h
RP2+931V8HGhjG4dwATl3NToS2hx0sQxjJd8+AZ5wXpEcApGMB23qlDB4e4gFWT7
5hyg1lGDHFZfxLMl428BD7nz1n2PVSMPfZZnOPUkbT6HmfQDoerg7XcSA8XNFb5O
ofcnptvf+jHkyt/zhUZ7sykTGSv/klN5h19X8lf7qWE2EP2fUL/jW0P0ZyOd1t06
S57VxiVLC7ZYhNpuAsNYzDllljyEc9sQwDC3Eg0GTIGMWi0r5++KYD3akQZllJ+j
awKXauruy9BAwIrRmMMN3uaAp4mSw+6Y1GMiN/fVQdDcd0c4pUUkRPzYu37Vtj6L
x+6c+ehD14De81QPa+HsbCP6Af43WoOeCTs7RixaclSPL1W8GTj5c1PaI6u82gH+
YQPc572yHXJZ+sHVA1KBFuwd6Wc8w66otMhrPFojc+Vtib/dDDM9kDEgBaQnKmsS
yxw0hMq9IRZBvhInwyDfgXoRoVCPu2g+SKb7DyvI1eYPuTz5ROcIhZ7s9PtafYZe
Ymvz69pAtUIoJbue9939urow27ifdBfgTGcCpffBbXrMzBjCbk/OSJ9e8Sd7UwEG
Avde2CPxAYGj3rja/KEAw8nt5K0/pNa8mYu5GIz3urwL+cZouhAUSt4bw7mogniz
HY9XWZwQCcG5CKKZ1mUcIKNuFAThTAEIGCcdotXEW6CG6NSpahKuU8pJDgtmF+Jz
ACg9SzaSh6IhjKD9PhbUxVWg1765vrgKtTRe5ESGJvtJiJn55E2J+qwwuAyx8V+4
OZaPxlLEmTVZMH7x/853v82H7NOcEHtgj5YTa+Wr8SFgr+blhHV9CZgrzgYakjKV
Gmr1iAf+lfTLpiMxg1P1ByM3yWkyylUgw6xee6WQbcpQT06iO2Uah+7vlncdnJm8
lkuyVyMKL5meqo5OWZFNi7zf1yAebIKuO6MAqv6UMxvbN9MDCG24fWUD7lW3yKkT
k3i+6T20X+rSqWnBpLNOtNuAAPSn7wfHd9DXePRjFg1rD0hUG8AwFawLfhYK4Qqn
dh3eO6SQXDU/c4QFH4CF8TZdZeKziuqgGpWNdIJ75wx0Zbm69WSY0UHnu+ZnL6s5
dgNDPr76qaWh2rAXUmibjwUSDily8jYDECXC9DA8P5UT2X99kwMKiiGCBVXaOTr6
MY+b9EfRcI6mdZhyVajGz0sR9jytUuVK377HG+XSs6bC6nOFgVnkV3EiKl4jqgLq
YrkN5p1DHj6m1C+BvxpZkQi3ueO5W63YK0ZMw4wpPMT8Clhtgpc3NMprEWPm2RAl
qdcXjT5ud0VBjDhH3NBImIdf1vU0kj5DoKbARmh74zPNgLRuz5RaVM0V5Jmh8JYX
840A3CsFvM6L3V6KLbENTAftLSixSp+KhjpMhSuQWBl80VIEpHW7X15KSAdu4qt2
kU/Gj+NZm8EGC5i/XLsEChZGriZrvbCo9V5YHhG/FEBBiMu2GZWJYR5erE8TpkzE
0vj91Cskt8f8bnMyL6kva9yN6aey5I9kU2Usuh+bvUA4N0x19M2G1No7rxPZwwNH
6hsS6KnomAQQxXtRy4OZW6y5cHKvfresDxvbkS/SNsQ12q3M7oAxAvHupkkYeuOA
qMmq+AaMqtqY032EVxXnZ1DNR4wgZzU7E78c99dqzL/FqhmZIIY5lUEtjLaAByFk
Lldg+rRLVwkAMEk/kyZWFVblSJEHY6hokGLT3Ik9/6OtVvEEwbsY5SuMHB7ppXkE
HQIS3Ys5/mqUz9WPp8QzGzoqov31ymxlOyhp6zx6AnAKcndiqOX/s950kErUneLy
DW4jlFv6AfDy/dD06Syerr9TCAJkGdYdUKWCtHFya1U1Rs+/r0/222F5SKGOEBzl
JWnFnsl9V+r+6gUGHy9YqCmwHuRo2dUT/ndtAaW1WJhWTZpSRaZpncw3w+RdDQS8
aPEox8PXeG2lK+UvBnEuc1QH24cvnpBFCWixL/eaT5gLaxeB1qzJQLQ5Lz+TKEIf
YN/kxD2nPaurtwxzhIuU0iMxX3F6pAxkvsagwpunN6Cbvby5VdYcyKYjHJy7AdNJ
9nfi8U9xuciAQCl5rUhftmkSc5WMFFZxdHRyWuHGnRIO5meW797ewV6547Tmk4YP
tnjWJkCdlx45x7W5BLCrGo/cW3Aa3HYr/0CiHjDqZBm9WUXR7BQqc69ZDQBg2gRn
Gg6fslaazVnX1Vp+55sBJ09rHXu8LKDXMoSziou965vqqYp9W1XxpZZUwCYscwO2
hAe+G5tuqKCXfP75WTtduO6dFbx8H/zg557wdxyRQZtIrl3IYK+/oUiU4CDv6XkV
E/CHEzepOy8sQugTHfFTAFws1KfAbc4q7ViKPFvhDBuqR/HAbHyvNMp3PpdQ845z
/LwuAO9+yAh+l7g6lCf23fCFqqgtC+glhMUHEvQrAvhD9OxxGBGg6e1C6ImaUhN6
2qaPPqj/FM6JIdEoKY1PAtNZvO/HxcU9Pkp/9hyLGdkdSXE26bGmP3U1WbPeZCuH
rK9/Jp8r3kACHO/1rW0dyrmEe0zBSIF53kakbafm+Y0aX0JfnJMXVyVuLPNXQPm1
T7f+F2NXd3DcQI8VOJXAXEcHt2++boGxfaqQvvvdRNSvQomtJJwFxAaRhQht6dek
ek9lrhO6splKcYyVlLsgvgLYBkvvz8W0GoxuSVrpI32kLScFh5V1Eb1pL7eIx91s
/7/PJe+5VVXD+dL2PPLj7Xq5N0hS3cDlaKAAPcerFSjhqXOFRnd5TNyEcxa+jrg3
u23FbnStHR494lmqc34OFxtk1nOi0/NKBfAvitSGPm7AZqbW0poPXWgRT75gyyHE
Ddy1TxDxU38Pc19LZyhU0UUhT21qOaJkT4weYUBr/nlgnkuIrh+0ThLlN1EmKN6W
UkfKvcvVG2AQzPPzNEwb7TZVnoUPD+fvJ3MK8I5w5QGHjeiSBHBt40uw0g9tU9CS
yVrxTam3mqi2YNnXGhun2SDdjPMNGezv33yjWK04p+3OLOy5sOtsXR+qnz2XqCcf
0ypPC/UAA4osnH4HrLy6ZxPl34ks9HtgQxwjresbitGWxBdawrM5zQFVGWwRhfm5
WJmg01icRmGEMRfInQ0X8N3P9LukWRfeg+ZSfo2fLVBFBXT0JThVqNuDYXWQmWf1
8cgCtDZZRgzhUDN+oUeNfdJGPaZFfTPN3KVHMMQioFVBB717yMyMD4cSaDxGuL0Z
BP3cKpHJ+ovubPnuc7uRnuzRx1lrsASMM96BuzBhspEwdXjvaW8qIB6dVPaCnkj1
nXdGbpAX/HG652uWXTJLvMONPr3tmYcG36v7d89stSizMikuYYP33GL8SwvV8w5W
MirOGfaLzQpVf92/+n9/RgdCmDuTwEXZjaHgreRZSvhztnnRQaroCsT14Wv7q83I
o0Pe9KWCDOii0/uxZqSiwZeB8uxW2Hfe5dsekCuv/Ot+QpcgJh6Gab/ybR3kZW/P
0o2m54hAgLPYR0S+dDu4nT84rlTXLLs4i/atDzDSUHwJG35CKBVaH/B6ym/WQ+HX
vPplTUbkDD/KokxrVSrLiD9J25IkSznMv1iz6ZQohG0+DsICHXZjsEp+QV1PFhfp
eSEBnIP+NbxNbVr2C5hUduDGckQ/qfwVXIwylmDBQAehWAfnYOmpR7cHk/ogbGN5
9qQ7+CB52SU5lQXG8TGBTGx79baOPHClqzJY5+5d+ccdbZXnSKIU28RzyUYxCKrN
ihg3P1Kj0zyTQJTPsTAI0iy2s7FHPgxLYP0yPoZTvefVGHKy5A368mQLtPbx/LQa
DWik2dJg1KGU9thVvcnGG2V6gpm+WTADrMELZaNg6m75gpgB6i7ah9MFNOvZjgEx
RAvHDmCCQ+ESw1ffUZ9QPQYO1HkYUU2Z2v7+LZWEM7mq73xsJMAUKIPR4AlZ9Y5M
f20Jnb7PIvjITJyNJJBXARWrucM7M7zd+WicH0EK1ncFw1e1p1xLbQU+JqW2IwWV
hfrHeYozUSQSi2zLiKTNKpP1FW/ZzGNEfY5zGtlGXlkOdRBPGoQ3xNPwZrtHnRB5
ydZIDdL3wBzIJsRbvzSvYKIzeV19WuqO+mWr8ytXlAJrCexL0mQFKastRs+o7vPW
H+qDt4K7xqQ92CrreGqp9bEtq9PBC+grIuxN+6cTkrIx1/oFf+f9DKGzH79haHFb
3xbfohSv/vtzD1dfZ6Sath0iEjJIp3UGb2I96I3qVoWKAHk+GNwnkZNKlk+wtBBr
i9xoKiX8ZExbK+sQPuS7DWVFgCRYHZ7BQnPKmDnO2nyl3fjz7rbTtOryw9aPlMXJ
JuJVVXo/vgG4RYmLhgXzBt3g4PDkYu+Z+lIeuW4P16DDijWfljF56LGmMo5mVIwW
aZ5qFohUAI8JMzsrUGqebBmw4DcFtqu1P2ZkNGXHSKlHURnxJqm1AydVVxuuAion
TI/JwBGki2gCULn6dIiYy5C1bROP1NMQbE60wsEwtvRgQRhb1cHP3CjZxfNzDwgt
9geZPpiVpXXZRTldGoCJwGNKuFCEUdvaXah/n4QXPu4ri5WqPuBoxsORWAew83il
evyylfwoNN6U8ZfFaGgWLuWI36JTfl/eP6uxvnZ1LcFm/mD+IND4JvvXudOgAyOK
bcH/iBAo8A1QfgK/GAXlqkGAOnCFxlvA9VG7UC0Uiyu1vfl7ZvrIKvtaKgTknQb1
xD52le4CqhKVVzsBAiwilpZf/6RlhZdrBS3VzF7GXbN73SruQLY0FHvM/KsOdJIa
I4ii+oPSyj1SRTpl3J9vJEyStM/9flLXb7tpeViKvxIv4ogBZiKMvc/fS+sSMwLf
cqKM7RRG0mI0j2BrpSk2KVaJOSSMZ0X+kzvwuXmICsDD2rhU810g/OvkDINDCn5l
Qp/xhDf5w1dzKreDMLUX8NWDa2AuTCiZsjUAJo5FG342MHKBBY+X9AX4EW1277gZ
rFAkuWwusTU3hrshZAWzWGCDAn1UM7C8i1lAXRgfWvwGoHToPGFCO+0+AI7Z3vZT
JgWJaA6BchxvJtmJkdNYFWuUwoLHpblTCucaeZCxjLNP/+3x0jlWUYz9dQplgYMp
eE3lFdjHLrkGR7jlpKdbOBnp+zqSmiKjKOb6frmgvVgct46nxyTduxVk3/WP7kdT
vk1BecpbfyvVf85FiLy/YCA1CCy55HHOxqc1N7HXJBFWRGLTa7JZ0VD11njbLgKB
X0wlJ+25pdlT7Kr0Tkp1Xg9wdc2nG1hjdK2+Ihau0WEjQ4F7CHqZKxeH69vqMykE
kVCiahkjA6Oa+zG/ubcIFBZG11g5o/YKPhZS0/V7gLKV8h4CeVcH/Tb7JSoW+iom
eKApSb99TizbGNvouTi3jCdP/l3qy731+1zgGqyrN11QCon80u/Qkq1ryzQKgacj
2se+bVNNNbyvNi+EWMN899JbykXXCuuQKZWc66h13VrI/HuxtZMQkQfbi5u6zrA+
YLoRvg4JdiKLoEcw/uT6Db88Z7Bfj8IEULWqUeNROKfzsdJxo/ARbNnNWSYBuePb
yTMtnjOhXPB2pNirMELE/wSak1+YfaV9tgwpdNn17iJhtmtlQGra+BjGqdZPjx6L
TUYmeIS87xMJOp1P1QKdrQ7Gy0OMliq2KOn2O8y9dbfm8nrZADi1s9h/y8jSC0FK
sdC3e4++5nxFAVZmGsa9QHLDVXJlKpZbQAgiu+q8mivG2FXwhSJM3fFe537Ak78E
z+Ah7LGBVEkxXD9ju79SXPXP2l+WF2ml2Y+Mqr3LQmCd5QR5dGN/G8JXku5/SxF0
ALV9p/kxdK4byLuChoE5JPoruGUYvbstpWQbvSciFKj5ZO5sYD3KjX5htLiptnAq
QLxxdQyQc1px7x8t4h8088rAwy5gTaMAWqXuJLOU+O93UrxERJZ1qLeG3mdAvr5h
DaGNV4ebqqFXTCYaQwd8oNcZk5dWNaiy3PESl0eehU9LRw0sx82QNEhDm7Dwl/pT
iutvWOqGhND9awiKfx+Uor/FrfpvoOqcRQUriMj+FSB0jfUnHAupNoTHtBWKAVzT
qYNN6dxkkjbRLUhd7MNq1GDP7Nhrdg1sPFS6rMpxai2QW7mVWC1DJ80mZz5V7EbA
43k3WhQtA6AlkSweTJBsUYV26+DqdJyIU4uqkskoWH0dDbpuxsbg1Prfk5ahmfPu
gxICg6zA/oc0s70tEmqfc9/xpyDvytgz3oGtKZdbXGJGWEFLCpG55hAelUNVmq+o
TzX692WpY22QON6HXwbblCsKyOKJv+QtlfOpmjNEVVDnk3mW7KnLtHadOCCus8Fw
lIgacvP8Wmc0DaerRbFpe7kT5Lg+cD7wy1EnBtJAOFF4PLCRY+0FttmvL3kIeNS0
nvB8ceLJTWJc4J6oMfeciOECjTlBsqazsA3bCvCms9Y5Sne6d2Ejswl2t40YLfnE
eFL+FcJgggLmzUilv19oV9caqyVsCVDNDvYxItQ3NtR4FNcNXrbXAutryU0at7pk
aDyoPPFwvMzGKOgDnvFPKVIqZoAeKNcmrLohppQ4XY57raJEll3oIBQgHwD5sNiV
1NmpIMH1m4B5O9Y+5SCUv4ydSj6tlcf7T8jddBeDOLYMStiNHIc3r2VA8Qxw71KS
i/VLvbmFUEINx+sQH+c+pj4noByG16RU6f9tBQTDS+c5i3VW5RLPE5a3YF8W+UkY
+iZgMEIrLBeCA53BmLujfkdJutftobDRnbp0W3FSGrrfRIA31Crmp/nPig1TIt1o
dvrh1+CPh941nRwAKdLP/rxATPsYltP3yJTiACnz5QJm6VeJpe7FGwIr3KtkvHSp
3ER5CqW+26YmikB3Q3ZPrpj+KcEKlUK5Bg/qprjeypj+bI8Rj20jt/AsWjBWyGu+
VepF0byU++PWTkZoyfE+rkJXkeLGRopPsgCbHWMu9nhqnFATj2eAS9alw4wWf+Y2
MN8x3cfbtW8pg/S33k2kixRVPllDenQYaURlwyKH+R/N9tXWHsslKyHtsu6TCkTB
gFI3FtePvy1jdKYr4cs+fyuoUI5ZgTfyxQUvpIasdO5qYA3Bj0ER4nQn+037U0Ce
CT7JgDKvPCwUwb+QsegJX+z40OTbsgdaRamdA9pmsTJmgT9pRvJVjHrYB1J4snGB
QlhpyZb9gPUGZErpJQWBLwa5ezNOuYCVnr97pBgdGk46jK14xa5Ga4RV2DfkT/IQ
8LCtqd6yOqFXCCfmtDtFpFd6mP/pYyHCEy7K8Y3l3+PsLQ2TkopK0+Y7ZM4Wq/uM
O/NyrdNksKSo+FYy+odanbTCe2txC7p0pQdZLDWac4KK00/xsM/7y7woepsp8+I4
6hv4kscOtPYXc0lbpDs++OcjwRVM787O/U5TmicuKbyIMDd7/b3iA8p+x9dordNP
jiA6AkORizoAWwWravpD4imoX+1t9iObySIUvnufdJ2pQI/fFO81WsRR/3pppIwT
Ol4+/8Wnt6RwTQlXOokrEIcuY/M34t4rNvaMienBHfyWWS89Gnwtuu0o2oUhvyp0
WeMSA/9VmFG0QSbCEDt+BB3njtl8CCyR+nt3ZGDEvPcrowDD7/r/SZciwYUioCf1
nRn3UO0/XpgOzbnFzZaPXPhaJepkD8Y1N24GgRPU/tFMi6/+CzsxOr+vmNdAu3r2
vZotKRGuydSOHT/EaG+eZNK14KjtbnE1x1CukkL8Sku/6zRaVq8DzfMw7sScNefL
UVHO5G7PGit5J9hKNL5ck1HkJO5osOtk18Q5FSr3VnE+b8Xl8lucSIhI+vIYLoTt
2duggmXTF0YPA4aoAksdTtgXVgLS8TFdD+MUU78f1t4GvIM03+OiTWgi6hL5+nCE
EwD/74ke+XdSSlJIJZXttSwwA9KWkvORNoQsd6XMImnGS/AUOzDNn7BXHebbigs+
itBPJ+srX0N6zZc96ZztSYJ9XtLLSypFIkXP0obIndN4PR5TBSA06IZRnESeKYGu
0hMcee4xuFjU7LxGdIQXkivqqUtSDI7FBvSDrvFrySNFbr3J91VAYHRmga6NBKlR
DsyiINF0UKDTckeP9loWD9EW1NFQ1A8AO1Z9D3pNWQlzbGSSY+4oJe7ixvf0aO20
jM1VUlm7C//GhDSzy6t3sOwFMswyBq7TJdqcnOvtHWP63U57tAJt/+t57nhWMOcc
gp2L8RZbzWdj+JullJEgjgQPsXw0gGqnwydPeiK31mz1ALEpcN1kbmJdD+2pNXmr
sbaFyInddsrCofqVWlKwNykpVTnWxHFsH2F0wz+WeBVZl3MFPzC5Pcl0NXdxSYdb
uAcqk2GTOLI9Yu7D+ZEbq7SqufttaeFLcrvSgTHkkTmdEL8wTJQM9SBy8cEHbY7Q
vl22a/EPttjGS+PAlUT96ltXUhWKXPiItkgvsGA5r85SVshoSlxDrE26245ORza+
yBmThzCPlguW6WgtmtA94hnlY0GFYUGJnqg3gdepR5rU4k5AVTxaPYZHOkslP5fn
t5kOdlmNlUDjb/a4bi9FUV8TjNHzRo6H2hzXccyMnVNC2uLF01j6OoLNum/u8PIL
f2vaIu3GHSUw1otOXj/m43U/Qj7nogQDy6EcArPpoHL/Naoic9QXOkEMWKIgju75
b4zHmetxiU12IkTIX6gDGK+8E1r9W+fKmEZGfNS3ePYvqRaU3Tn9do5KWvhO0ec1
Hwa3e4cLkz2KlbDT+xHmF9IxKY+9roY+ZRTwqT0/8N7IgI5j5RIDiixRdevj6EMH
tc3hvnQ/35v7m+7qp8UvimVPv3IpFiX8Tlxslq5dkXNi8tQrrK05Zx9Zk3lddh3y
Ana4e4sr8UL2kv+l0FIdIN5qQ2fRqmslqpi37iVyhiLIUrww0PJsORdYVwGrwRYK
QtlIE5q/AG5T+Bo965eU3f/9AEiNuSasmz7eBdX2i7xogAXqkRZTUm/8vu0XOy5e
4SviyWJ8Bgnfg/m22OwnKLP3tgf6PqKsVPrKk2BFd6CJJTuT/vhvjk/c44B2EK0a
b2ZpZ8LKe7Pmh5jyCm3Ii6im+cMjxrxkCmNoAFKFlA9ceyjEAgaQBCbQi3Z7V3SV
j8FV9WAMWLJCMfd95UBQAVeyKC4s3euMtc+qx+bFwB0v4SvYumegQWBABtYMuA9B
nNQAt//HulJEWM16Y+RiH1KyG4GiYgsPfJBkYVj/+u4zPHsjUjhxuS8V5qc/5y8G
gXv7eyOwk4uMbfa/I41hjbYhf3Hf89TLKBsz7rWYHNKqAN7rBo1mHzUo8+mX3ShX
fLinD3iZ3LhW6px7GY89Ktkn/Nf0k5SRMKztccdiG4jCmSkEMKaOVqXbSfL9PxN7
ma4wQdVM960GIel6TL+5fSBNnk4mAbDF2ru+PcH1z/j13FKdx4DStMNZA+DqzwNI
sTo5nxSUF6ytMqEwm7r80ABozQwt63K9Wj6Yd6NojtOmoR8YrJVz2D/2sshn8afY
2osQRCeBI4VpVWYHokRLfKCNEeCFKRdfLBy2QJIS6Cm6Sxg2cyOdnIZLsclsWh3l
rUfqakfuts4M5DGTZ9XWX84RCMSfdy0ruDAsYHP/wtXGnOGsnVbs4naSUXBQBo5V
ISZX+d8GocYdjGqN3U/wskRXmi0lZV1D9lrVBtK/+lqijMhBj7fmfiOpSPKcmrxN
IEcfOWKLosysK6A6hE0AP+CljUVmalPe0nOFWvLcp+cQOhCmvmHtoRDnhNVicRFF
gQZ0kHD7/O4FXTV2Tcicp8yIub+CxPtTTkqTHIFNrJPvzI34B/4untV279jy2iXq
LToheTB/f1+omEgmJ8RrFOBuNgIJmxjkplrMS127yab8O6hq65CHQ1FhVvQXwT6E
ws4ubCR/cPN6SAKpbPcgd3dlIOG8qRfgjmjk4PcOa7rDpwyPdxM7mkar/TBnfVte
EeIV3YFibuLCf2bkV+fKMZteB/F5XDH0T5fT4gqxLT1BL1/G/gx0sxpX1lT7CM1a
nRLpjfdzWeQVf7oTDkie7EZm1NaCDt0hp1tJg7QcLuJF6XvZqd7nDjqAiSw8wWfO
knBUPsTafWWqApoX7RIbPcocBcabVgbPAq0AXnU3QPnq8HTd+M0F5RlfNvRyS4Wg
uDWUsWcX5BFk9AF7Jc1d8WmiByVtbbz9FVWPBIhnMtcmM0TaDvq7T9M/Xfx/AGGs
GVbICx/0HaS3xNtBTOqZFFhE5UGG2zOJMwdPKcra09f2YkmZUNvWgj5uzRkTQP9D
NT6biOa5K04Stc6X3GsS5wtir+P9kNdw85O3mcTPbbiykDR6xjD92aTEkTrwNnNf
Sn0Be+2tvHyndq8/F3IJOMN5CPk3oRh2arG76JpLFJaynxEOS65ntgCnOHb+9eSQ
eM3D2H0LadE9+M16/duJrXZqbmwP9bvuEXmIoyJqfRvHScTcN88HqbA4SFPnoXFV
vY1QJp+F/1/QCnBVCUhaawbaWpfF2dGkM4oJvktloZWdS1U+CqKSzIssclyhvne/
h8u85mk/Qu/sJF7YiV95sJDIaVvR+OqOX54EnbFU4nZfSqc5ZZATeDC2N0dt2Djk
HBnKV1DV/p4vmsHWCr/wy0AzPSeYdKbvIwHkSHvXzQH4J5BzOWdJ0owEQd6od+ce
pVvOWOTj91858UZov2krHpUGFc1RDFdizkUfuJ9eA5Y3aSKtWmtynH16H0G5aoni
lA9RnWuUWpx2X8Ia9P2FtxlLdTCxzu4qj/ML/jXWeHL0vaHfCR9D2zj8ObaDEx8R
G3FZDC/xa6B1ltZhp7eUxpYmgjwUeAUNbcDWfsxP93yOg2KMMukVsUETl7R65Xvy
E+Ozyvklq5jwYIUOhz66OtDUaWKYIAKFfQNoo0f+HApHNGXCHx97/Q2vnvN8PKdy
mKdSMpc1rKGpvXrc5pXHaWZ4ATJMBGwdLaJfJEFJwtuNOwUedre8ip6VM6yT4vLs
0zCjz0vZ720Jt5auDXEJJE2Rp9+RckuvQuJIVCGbY3t0Py6LpVxZDw9r18LE8NxM
up3cY8k4XfgRQIBvfRfzaN3Gq58qBnwQexM6imQjO5GdvfkbZP/JccG1HMqP2Chj
Awx/Bb3n5aInRJayu2g8RWiPzKAQeJC8S6DbHs9PUcV7iCAEF8qACLRXsdYqXGNT
HrNdO9WLUwItMvdeEfHKJuAFlfuI8NoOBPTzMhUxHDhMl+etn9B3//lgKY0bwVt6
zSccrYBT2DipTql2F5vTEqse2gfuJ/9Nc0WDa7Td2EaE4rfSOAfV100ibHDfPax7
cpCclgXRrcyTiKmF5ep4oB+fCjRvXXtahUlRJi/8In3eB8XhvVFGsGbdJ/ly8nd4
wyBOHg/Z7DAOOVvR3vdlzIL2tJ6moFpNUBejzX8Vd6qUVFMYA2chNXSpQRpizB2P
3btTviXieX1OJkffLBr9HKnRskE8Z78qDoimfNro3OxPKw+TvKScP2v68s/l2GHR
b1Y7ndCTrvfY+JEJhtiu++Ig+Knb5iKqX+n+O0nWAQW0UFwyn8J7WxnqrAuYXZgZ
hMImlsMbkUPhaXgVYVYN+GbZw6Pj6zxSsBnbiZPOpHqG1pFExMky9B7fEksnbXoW
zJJ5Kl2EDoKfyYMTFS1ALwdU9qFFOyXG85lHqBkCDqozTclwc93MJfc2WhV0P/DZ
whxwqNg/tIUiegN1T8RBJQe4czsNh567mpKEkp/CkT84wCJqqZ4H0Xa93xcFMl+O
Jq95ec+9/jEdF6odcPrEDC+jyzXrXq8V8hal/fJobO5eOzlrduA75qigxB1VBiXm
fDF0OMJOMfCDWmBqVu4IiEckniJ8EqKRd0c3KrjPB1BKBWoztQRcij9ZLr44oPKR
9EGr3mHQcWt3IUx8gV+bxoWskOaiy8C7yrqt9iAFP3cQlXwqUUkHDyLzyAlqspo5
4QkYoSPXaoWo6p5Wi53X3aq6JYDjDG3UEui0z6cAvh4RwOYGIn+3+GqLuzr3Dme/
bTvEMPbxmLqtW5dSxzU4CYfJmXlQa02O3pHSBHeFzb4JaLuzNP/eX3DEIKcwTiGu
ThFksQCcdTgA7TZFQ3INHnFLRIhLubZLlnHQZit86zPs510FetCF4Srnnnd34nvt
VvNWDdvpzpLP5Yiy7xT+ZGgU45TPVz9KhhLc30CbAWb5d9T6Hku7pfY5+FVxxhkh
/+3f3tKS/srlFAQl0Y4jVX5JGJO0cWUXDgIdwQh7I54/j8Zd7Ba636ND8WKGTz3e
6dYSkb6Cvcxgko/61Yz1Vm64k/ACEUYqVO/QofxaNUn9k9ghxVv9br8fwRApZBht
+xV1khUqdV6oTnTUnEV5ZTTbwCBmTOz8IM5ZmionVdHi1+93+oaaKDHWHKPKAKfq
xqWS8GKvQxS7ezM7FmqZI0nJkntpCJSc93QljFgfaFJg0+Vpw9mMy0R8W97/rx66
ttx9M7IEqkavy80kymDBqerv+W51GtXfRIYgWU+sBl6d9ojRd0vCS6tAHfBX6EzV
tXQd4B8PQy3Shn/+NsXRfKnEtyEy4Vi1f8vvzaInKFToXDjYA7v07WNZ8Ny2C8SJ
/wT2ddUZVPKXYVnz2w0afuXeEhrbFxbXnO4+hykpVTWfrtcPe+Xj4SgGuCB4XrjR
n1rvseLxkj6AG9lPIXWqELUrPKYUWOM51hHJvs7v6OG7hwczbRNLh/OvNPCD9yxX
3cUrTMi69MTZk707OZPGgb27eZwrpNqpOcidHrLMW9zQFug/ESwEuuW0tzfiknHU
39q0VEV1+L11fX3uY0mG02mxkGe1cJ6egRZGE6Qegrq6RxrSB41AcuSsImkTZhuT
+PTpWgLADQLYPpzK4sH8AA+a9xt9EHbu3wfqnh0rtDNrsqh4r3mfwfK09+PC0RGz
h9fQbEVXsgd7lx880WmA/YyKAEVYGkDyijbelo1gHDzhb5gbTV/ZOE8mX7mjnWbg
4bS9tqcnVw7tmRbnJZY22+7a3pMHw8eUqIY5PKybKQj9UJ6xWXyZ3PSd8dElYKzX
vc1m4Qj9Fk5lN1f1iKrUsCvJ+TccMItYgroAQLRqYYLqEbHpQHWT578ZNNv5qmI+
MBnHza7pTfjnnCpU5PfR0N8PsgzCMaI+5C9NMjReU0Gx9miDfLsRpuCI1DQDagnV
g/QORIxhGSpP49hpbWxf1rSEFUfcKrclRZVUmSU/0MXfagTcyoP96AodkNupzCTV
mFNiYMwCaknVPApVJgYGmlxft8A0WdyzK6L+y6JR923GnLUa9LmLFUhHT61azo91
JugrqBj6WWj5WGnHa7XWYxXJ2XBr056VMBZ5/Y8zzR4rKgdIEVC2JWMJk4Box2ij
sN50hmk6o8g5H3Gf6CTvRdpFSOP8c8zATPIqo1i/WFtbriBFA81PoaeS+Ktszf+b
AbBS1wRzM4jZAE8keWwpnqkTaHLRVXkI6XpqcWNiYv2B9teI4z1Hi99sYc1KXWW1
rc2+H2qJhE6bjT0GCsbhBH8miitAOYrB7fmA+GD3bWcEOfYDMoZ+WAgcuAt4Fg0P
M4sx408sZ2MTB3tQTDicoAx2shGbAmGsA0WsPPRM8Aug68vFmyDMqbxqLvmXrcWL
E1QmJM/tvukM14rMwx/pjG2F9TkBNeLq7eIsYS8DlS0CCQHdrW6Fx0qSCJ1trEpq
jcckYFN8hhwDNvK9oObjpO4VScVYRZ0SmzM9gacK+FK5fdod0gBLqanubMjjtKCS
C5Xx+mywvVL/f5DDR0x2zgYxH/ecGKemlSUwMtj2S7hBkATJd324kIlxnduNP0yP
M5EU88u4CsQiqoXoPNwDBC6+DLTI8TBjk6V8jCYOMNoUZY0rz4lROOXVCUp5p++j
4iDH43/joV61+DnOG2bkJTOt9ZnZ6oGhA/i9CUYvFR3d9JZ6BsnSwv6SUmh7Eomv
aHqxR4klurB/uEPqB03ktrOecEuAR8RJclYHG/ygA78x8FTpUdiHoiIm4NFRA/CR
o63x3LFDgUDgkDz2H/pkdoDCsH6Os7rTGuXKoe6E/NB9VXK2+ICoiYB8IR3C444g
wHuACR3TFfdbjq2gC1XdIUKQNz+6qeQlrvsBDaFKOv3JHIlKTgPDM6cYWgeqrfzZ
IGpTtx+cWHN4+GxKuIqXctYGGv/wGDIHiWB+uMwQPJF7DDz1j1VIDPcdeajZ4vTZ
yyXmxEtk7xVQpvbNLm7xdhV9vlf1LTguWlYzOQwd5HqaPezrZjDvI2RQf8B0xwjg
nDPNJC5hgHlz8oM9KnZgWyY0yfQpD1IOYCiEcY7CnhP72ywFD7HYfiwjtgLqqtAx
9LaibBmLlFeTsrfBXLNJh0knoP9hzQiJ/CVNooImKX0sW4arRDkCcFcaW5GDFC0I
3lKU0fOH/yBwfMIBsupy8W0A4DKnloRMK4uDepX/DVrtlXXKFcxx9y1uaRXyaiDe
oi7l8el523Amdj/678xNNDvWeNYSnDyiJ4LyUbYjiYbwakVJ2dCciWYq0cZg1r+a
BufAtv6GAnOalkdV/JDdWtz9AvJsjBa8ji8SIIE0nUC7PyRLTes0rsDRuKVJvdhf
wzUrySYRTsFAbmBrDsSLbB+XAz9u+dmJiOyio4zTwlUJeZyDb89Lf0uDz6CCoXW3
j2s7mcJTG4afIDwfCSuYKPJEMOpB14PPQjGk/chMlrVasYuNpacygKtupb63EibP
bLdVdYZuBv5e0RNcEpfTQ/AGlBhX/cU8/We4QtveyYSjoqXKIqwZd3+/rVKQcW1D
PWRQ5XJ+KcpjzWgOno69soUpKwNFRMJVfrJ/zZ/DxHEkymE5tqHgo6hFIZE0lmNQ
ZLDNaKs7CG8bMq+qERnqdaSSjXUWB2LVhnbRdBpn1aWrjK2SwdjLgOBa50Tf7UfC
RFv0r2B814DanXGF47XiJ5BxKAYq4ovWBJK9UF6zESpWmya9FSsOCz1fT/LrJhoE
75uOG0P4/12BOM5EjEqdEh5Awj12e4O2nvRjilGgmm6jZf3iKmbfmtYbcEESuq7q
+J/kUMN7bZ8Aby6uQ7hz/emzz6FFsikfuDQ+TPhd0JVNLYoXrRv87wPtH5AeiOu9
x3fd1L81w1Mkh+81ymSvwdgXXMZU80o0RdsoTP+d9INzoZDeEmy2XAmcFJvLfF7T
JlUKTA43tyJrAFaTsg8G+bFUFZo4sv3ooHKxl23pxV++ZtIv13E2PKcp6ZZvXmCF
RwGT/ce4ndv83E3a5ocft3KMYxE3RBWvmM/sFbVzi9NLqkigCWyJg6CFOy1cAjZe
c8Un1BTezOL67r5RhY4Me6kFq7iZQ/cbKtGWuwh5njOXnzlgnNa/B8inu5cnq/Ho
jyp7jk2w2RZlUawDaH34J0zcUc5r8aPdCyerhHSOECfGrvzLrNevC28ojyisZouo
oy6EDyWdJn8S0yTK6i7mJ8u+2ZbsU0qt+5wQV83WGDRlqjXlJbtg/Ltw77QB5rnh
r8sqNoHExhmyYMMblDFBHkLA7MMPs8VaOlbr+v3YLoOguX2SqaceTNMZfqiu/bps
1UmwcglIriMy5K83pkL2+TmwwykPo8HSldeVkMTXUmG28rSLUo4b3mr7HC9iqTwZ
MtoIHKmvWLRN9rSW9DHv28lM7SiSe1xv6m00BJJgmJyj9Dq3O73FK/0k+IejW0Zf
r4oioa4lK1AupejFM9/hXJxynPM80NTvprloWeWld9YlIK/hXBB9Rf580+OylfF+
jW7bzWEqdH6AKYd0AcTxhUZTJ31oEg1wEYOA5A84CaIzMmeo+xnESqivMQlBqvOB
fv+wCKLm+HZeOjXoDhAjY4r5I9y8/IKOuh2Up8JcdALtnkiaHeNMR5wkiMbEd5CJ
chF1N+WQNwv8ERxHlKbwBDIYzna3it5/tlvDZd5L1pEHAiGfTxwsoDwJdeLxuhB8
x+9linBoGE56sCKe85PK2ikcvfWB1Xvi8z1t+HhdEs+Lnqq5QN9cp3Y8UIk+28TX
UePWz70lslZ/PDdEnZ6MSWMnJPHt+h9PHOgMpc887LisktpK6REyInY9l8+QPSXy
Xix3x453YRcHgqYIJFSamee8D4WmGf1ohykesGEdbQSTLdU4o8lLF9eOF0L1LbGX
qJEgP2iOvTbbTsk3aPtRfqHYATaHvQkP8FBXX5KAGn8OfMyPZX21uPI6LIABRidQ
n6SavRFqBYFRYmA1cePC+HPpuWGygU6icvtHKb1E2m0XXjoVoT1fY4Eat9BxsbuP
S4FHxB2iIXstpQgIhLZmOPEQfM6TRj1yJSl3uZzi1vof0kBeTUMrl7qmjd6t/h8V
jUJMZqBxL4j362eKdE2Fr5mqwwPUZC1TrT8487dnXVRdYcqNnWzr2/vYfD1oD9SC
KXkaBvwP+l5o0MiH1um7W4k7BLJ1QboS714DnD0sZh9Q4l2IJwdrZiDwnHDgJO1s
lIscORCOi4uyqMxd/ZelxersoggfpBfNfBEHp2R+qvaHYPvZuGZpt1lO7M4PKpp3
6jltXzP70MBdUfnAluY5aYvwZ4wcj4h9iwCtGyvhimk6c5pDGhsG2+MWEy+o+RJX
3b4d9NtVV22RqugEsI2KWyaLi/i2GyRid6JDO9BcUl9w3kNKNmBtotmJZfsHZmen
wG56V6FxWwH3Rf9wDt3EUjOLru/lR7fgk7NW0QIPxnaUA5CCWoX4q2nnDZiPbp+L
srqJCARopfz3f8rI9BJ7WS094KzSxmtRnCSRRsVxO14NtTCux0507KojYqmUniIy
dGq4rIbv0l7Ahx7RNPkwE6TYRv2TAMopHpByKV3Wyx3JoeDlRyMCz5NN/0UU0pbb
GS84Swk96IgZpKgfk24y5DyPr4ANPUjqKDiUJTsitGpIwPk20xBwWIvD9oHJDZKx
XzacZBjgqY29CevpFzLogP10LLZGqHx+cXJKyLpGlyLDC3w0RVJrAuladZk5vgcZ
37z+Lqt4+IjlGhFICOi6ALRPmgEisgAfeSgZeM0oslQZYQJ7yAsxULDYO/c+tmhg
VV1MmZZtNuDZBFlU7LFmv29u1nVSyrd/abRcRHERw2/Sn2C8IBJxJsWJlS5w4Lk4
kMyeg7GQizhqrxFSup6vPWpdKKJNw410Uaos59gENWJMcyi1C7WTzRP4ndPgiGI8
eeoc626A0+I9LiXrKB/3YWkmyBW17FKIu/EPrTvJu0DAYsAo2pfuL1nYOd+G+S1u
htxtSKNByAqO3sB+V4smRd2c8iveAM/FMx5oydqL0sIcqba+lsy4Pc9gu/iaSeoc
miRsU+N39A4YvVYLlqcnei1VqMjw/PKIbI6VaIT14fqCUNxHuZ94fQeB+/++WoEb
8+emqURUhgTqmBTDWDFKEeYl7AvzwLp3qG1tDjlBwmmZRBhhu4WcyKu32VbAgIBN
/tIJq7IsbvNtDTwFR0xX8lz8uq/Lio5tX/InzX9XsuLgNBjb0ti69qvPoeVxjehu
UjEt8lvOnj+RFD8ZcBTejD0Y8wqkPRC3D2+l8u3ZT+ktHT3hVoLF5QknjH/cLeTa
ULURqgQG/AwZhteXFQSuVAy8Mmw0L0G4BSxlYXcs9MAxAMf0NXqSmMxwKPdWxtV7
Vkhubw8hWGKeCZhSypvI6raFnHq7DJvNJcywzCFuXu5+CEUMCtSe92tLXCECxGbD
gr6G3hz1ppWW0w16YCUcW0MugkeTswXqsZmmkfMOWUwSuxaeKq7UZxGeKQ8M7nc5
iXE+oRRPgMzueQ9qQKwZFmeIZxHjvzzom4td61iHZHAeJ+Ska7QeMXPF9Y3k7vBK
8QsIrd6BF4O8c1YpWQGJECgAV+m0Rv0qqsf/0neQVLJg8aHzkIKMo31GnZsAoEk6
tH/BuS9ht2xTGXDaNqNG8sHqMedM8imC2ncLYRKICKyVXtqVZ4vBIWR8a+A7P22W
U5WoQXypEa20YEWiAJdhAdEmLT0fcoesIoeFJdlqjO95BqwOREHa0pS26WRTN1SD
jphrNhXztR1XS4kZyFRyhyPtFs8HHPeGthE6zAt/bDuc9egf+IUJ9FvCBNy2StqO
Oxc6idX3vkBeNsoVUCD0R7A/xlowLW4w79bZGE/Lcx7BPehXrXJUAmbdfhoqVU9S
9qxgmHmkZ00oZxRw/wPSVY/k2fd4Rlv11WaumZ0HI6jonZaj6KdgvklqnsQMCapb
LEQ6HRJmm4WcPYLT5jWS5iCGIg70fFGiBRGovJcIrW6F8Wd+RYddxlhic/5CsluW
yBVeejx3BmjvcyhytAdimffolsW9mtE0D43vfq0NNajkAVqcAuNabcFLiwKJr5pP
/6J7Zfa6m8f9u/YgNzueWH4ArvzSaQa9lF1QjfJ2Bu5F1qahhEFy6ccePBZT1+e3
ItNI2I71fODQM3CGrjLSH9pjQNLQlhDz4+4ONr4Pp6xJzR33hXoaQAchmaqI0dZ2
3E1tTmtSJpiit6fi9VsudopfQLaA9aGpCemI38KvLsHmOsDT7KZbP7I03e8ilqBm
ietizNpHinxgLKO/O+t/46TvNGHQBUoxcVKqVsm/QrHM+fdNiMyfO3pv4Zs2Kimn
S35+8mVbOIEJfS86DGRRe2bgSzW2PCHmrkeDhuoxm2Ow61Z5vcWULnqzgpo0XK8w
yToAigTwfDVidcBC2Vc5RZEO8Hxob2r/xz3rzZowdD9YWV75AOjZMhQihJtwphUg
sz1Jd1nwwCzZYqlUP7VZQJNpTIHrWp0gJ/mAcNM3BdVQ4O+Fb/9DWYMR907cZeji
00z3n6kFUCMNY8aacrzuIXpkGIBJJaLKa2ukS7Bj3OQ0SuL9UiwU8/K3sh3+uMi7
KtjfKQn9oo6WDh8Y4vq3/DMP/n2urXvPdvWUYTiS+WrJyGeTfck7UUHmuy4Dr/Gs
IePKpjsMwhA7tpNKl/JMLW6X4+ckaonU9K5gk8duGD3cSyGukYEU9MFZRlULSNsH
/k/o7J+6LyrvtPCtDdoXeXc9DJj4/T1n+EOV8UCP6k03VOvc0oxsXhtvrgAI7CrZ
dTvRTgFJb/gekF+qHDQcfQMNV4M6uECzSVJgfZEjb7Bg0jGfUpQuEx/7p1DbzLpA
1ntAcuKWuZhZ9vKPbEwCzWWiQw1NWDXU7lKVNRwzmak9jso54gsGvNkIOpEzoNKd
xy82pWo6d3qjBcLCKXlWnzQWQhrhpjpTgyDlE0QW+iLaji0G9D9OwWYV9I27B9Y0
jNKrkI7JAvAmG2HVRo+1j/K3DFhDn3S2AOZjA5E+Uw+jzUyPEcJyl8yRSwFJI/Km
4RRshQBpB3OsOn6Mv6Z5PMJo1667qcyE8J9fDnvNKeJ92DDqklRewiX7YUFgiR0i
iqyC1yrnbPLOixBpSZxLBxGLCWL5Gri11pYR3Nu5zyM0LfmIstHtGY19oPt4J1Tr
dFCZQiQ3s5KRwT+oTQHedsaripnz1kL8FIpPb1806N9c6JxM9kMbqmEfSafsUA8i
F+KpPvFOJ8Qw7FnXHcRfqQMjyGQtayM7naZtIKpDBwSb2otryGyMhP8x8S05MD39
c5F84js0YW2GOT/7KHDXwZpzjTUV+2YuBcUR4NMqyqkKzr8SdBBDjC/5CkoQzSZu
8kiIJM535LjtZah4ik/nkVfx6lmI+wg/EOrAb+Fl9NjOeLMfRdlCqMC0cVJcP1DU
rcMff5ifCznrq7FCB4jOaFI2E2a248ZL0SAO1A4eLkWeEMbl34XcP7Vgs6bhI7Nu
oqkJja/d4vgn20S8nGQU6VwfyLUMZUdOc+nX4odBAjLJH+eVZ01VTuwHlAjlpgvL
IP4aSwOyr1/Fjsup3fQke7btRiPqXoiWHWr9IZVNV0gcCCro43Hf2AX4a3Uzby4+
qpctKHMTIkR+5Q2LbnoOhGVwQ8xXNBWoPxq5aIeGM8LJp7OgPmGrS+HB+saGgko4
BBMVSpG1tHPdQv4PQwMIsvBfPVhhM1l15cZt5vEfoZ+2aECa05vc4uA0Q6t2VHAS
AMhQD2vRhqtUIk+DEmRC0EULOKbJOm298pK5XQS0qwo0NQ4yR/QinKnRaxCVuEtj
au/fBncW/E4dJN8M3TtfptUkF9v4AZoztW066br8haMYaI0Qk5Cm5WR4+4jK9Ao6
rDyQI1FkEkuQmt8o7JvdTJz7ACtI/vcQ4+jJuMnZ2QRyGufPxk4X5XgJp+3UwYKD
gYrD5ffW+WQ71tzvMiIYfaHLaH5CWpwmgArz0Q4qmmChdK7+PWf4y0lDEn06jb2R
cuLfHFCr6uk58HnfaKKd4rVkwAYY5Xoag8lYJolgUGX6aC/iUKuLzU+hcyh6taSA
FvUWhbDfjEttQ7sQkYF17723v3yaCpHHpTXsNknuNl93jEA2W/CF2BDry4aUCQla
7Y5aqBaztHiS0iZqrIYuvT32x3ScCoZwaFXKidfBHEluq4JQRHs1WbzBtXJa3thl
6tdu2wqfclBe3Z0qAQNIry2Qb9VxiL9axiHG+ENgf1e9KaHWWq5JTp/TrHu+7VSf
Tvp3Mp0lP1pyPiVzE9Qkd2tGVchCtVKUvJzkQsBtU/fnqEuwmSwEAfKpWpBsHZLV
RHtFbTpq/fhfpT8YAVVMrg44w9Ln0BccXy4C5romISBmxwdaSvGnSByEfcL7q2ma
YttMWYfYWxQxM6OQw6bta6Go08cHL2udvAi/fZplAXVmGvvVnqPwH7PRLDxLhU3t
UWXYBL+2bQ06KPvw+1nnVRWT+k+T7UcX6e5oKrZ6Bz+CqkPOEYMoyyluxOHyEzto
7CakwrEH/NYcrgk7AhhGJ53QpMFKLeWaTKSpuyJsxUi1A8QfVJSARPyOw3TheyWC
MeLIhaDiW2/dLr44fWo7uK44F6/EkeZhEh53F5q01ldDBc9ODacsWZUnaIHnqFy1
RzyvrW0/uQXmvbms32/dE5ZvY7W2JiEQty9+xx2GORwGywpJk10K2YG6NonqkxZ3
WCmcYq7ZDEBhBxWEiuy0WN9fbmBc7Z5eGZmNTczbKJTlXV3CiytQDcoveK3rOtfo
Ed7ckIday1YM8IJ8hOBzvd49a7k/9OnMsz9bR5xhKwQbyJ8JOIEl/8wU2D+9HbX7
3nRlkjugmoaT85NgzhNvxNkJqxqE+qBGlqxjzRJaZqPyS+46Q5JwqNbG+lec4WA8
dCe5j2077b4Uf++3/L/EOIdpA3JCVV8SlypEXIV7xOb4xHGYUhFgzRFRgQuhWxHt
4CgFYXqYf71dEsa7ozhZogFbmeRb6uEUwTCid12HJPB0ss6YJh6ci0hRkf67sv12
idyJRbsdaAkQ+pGt30hkmtzS9uskMnK6NJYQ1OmDYPXswQBtLWV+kvL1hWf3PgHv
oLiUuH273WW6SHWEqMFw5aT13vHGamTOqlB68vlyOy735Ct6F3BPf8nSiv/s5at1
/u980rcbd+IK+DD/EE3+O7QcGPMy10P93N5bme5Kgrej3jxrjXy2QbDyVwozR3HY
l6oCnthcxzyf/w+lQ4dgKCZS1a0HQ6oqbGVKUt4Af2ZNZu/wh1IRrC06PmNJAF+F
GS1M4N3c+6rh1z5EYHnB5nAPm7P2NSy5IzvgarGwE2CqXZ4bPKKM0NySYDacu39v
NYLkrZSDuVoOsWtSCWroEYtWtjH8I2qNyatej2sJ1bvBSjpEiNJZTsfH6k0nzd5+
NY39J0srxr8KoAZMvouyFcsg0YIr356mu/Af5ijISWXNYmfgxQuxmy07AITC01K8
YWsMqhmHvzMO9foimRWV9jzz6iTwEl8JuqT3SgN8VGxhPljg0ApzSAOnTH5KGdZO
3C0soG0tWY4J/TgsO+fgxrBp9rJZKfKA/UuqRWdQo7qCDrZk+yRcPuoQCmaf7j6q
BcnMOc0J2x+gXlVA5B8I6T8Mtq9nVD5D9qqLKxFFBeQPWiDp4Sg1eJOBVuIHfnHg
iedF3Mz/g4vJ51SGztlt8U5ci8bLAcWaqrjcv24kDjJvCOGG8QSRFEtTDGpKPqzW
599+oQCOCquJVCDG/JI2tvuJlydHGhqU6mjwb+C/zAmEUXKREiT8jrNPbAmsn4Z0
DUoMgSD8dOSuvqjBN4CZri3Xf+I19pki2m/fp2L2vSY84atZ+scxLV6mVLKb7grQ
XD5yX2uRfwaoh42HKghJosLUqBKOeoHRRHLfSpSyJxyxzD4znmY/C5Feq1qIk9R+
4qCtbcvqO4hdS6HFdrb7z6VOvrlHU85sPhdvqNQpumZnjBiZGgvh4CAsx2kFs9en
ECTCzNJu3iw3/3YxMN015XtgN6tuoYD8GjOxAcMv4w7GCxVlqLfyMz2kgFBvoRed
PVPkxPFWxnFQcJ06VO8pTXgdqEgIx8otWOGmz9d4V/bBss5nU/OTrDF2VH0F+4dD
lV5WYITzgT60jGzu9Sdtvoxd58x+h1wmpdGhAKBLKuJ4ZtqncBQsyVWzNysLhSXL
W25Wf7Loyavk8sD4YhD0jIgx/1RzMo9OVbp8KZmo0Fg4zaSJVmivA5qSeu2aIpLO
pIsGpv0GE7Qj5AQBfq9qp6JyEcfq6aBGPyOIGIzMUakiTVNcoTV9SjbvET1Blth3
G7cxHzm/FMVJ+ZnwqbsmSVdWyq1eQMFMRkp7dBwUKKHAua+VjAq/tl6zm7cOKGwo
bsq1CtEQJETgQdWI+Rw7Xsyq6TJklKNIrL1Kt+EWOkjBxi9QlxFtSQlEM/4N0XDN
l+Bo2E12UtfMWXPgBCNPbldweyy4s2SN7Uwbciyd+FLcOMmsmXfaLycLz1tV+ryb
FZir2qUuxwBgUl3COsVDFiWl/WbDMNg0QAGesvGYvnfDPENHtdUVror2dmxiUM94
9zhqjTPUzoFs2QbHP+KKCUocv8Epx5VVHVN4MqF0zk1n8JA+E4gEROKd6sjFBJfD
kJrdhd66Sbs6r4NWETMWslAkEWf/X6hK1dL5xmDdn+mXUAFTaCPskVKRZCWsWws6
vjvC6/A4ilaQAjji+vUgd9dTKA4IJfokqwU2rULqhFrqJuASC3fhncGHpHIPztO5
cDXX02No7ZQUdwSNOZRkNtBsEurtzRarW+2aPWcYKJUeeujHi04j6/qSK+WCCCjq
H9gUkcucuoA4Mqt+LlyVZSPQy6XilU6xZrmHuSPAIBfOY8QqlaYsogdyPkjU2xcj
NNYD17He+4koRyed0DnVZFly41qK0nLxLPyR94c+N12oLBI2kOboCR4BmixbDmo6
7o13mlrxClyuULxn4efjs/BD4lyTbDRPE+5Sd1MNedy4HRxHfA15D9g6U7p2hVCq
BcIZLsJB/rS7vm3ZD5RkXTUqLUEjP8xTgF5dQtVECYb3wNdQLpdRk1Z5zB8Ouy9G
aArU+cgru3Ze0FxK+yuEIeE4cwSOjwFytDmNqQDsuiac6s4+jpDG+FxF2ttLS7kD
OYCl9eYL99NGB3xSlI/fIkayv0FhPYuP68I+ZTRqCyTOKpvFm/kO5dmmEC3JifvV
MSJJfZdgeWItlrozALhl70RWlIcynM9TVCh10OEgHg9tPyQZSHLMTq0yL8qb0bf8
3uDPyYsnLr3gzouP2Yd9jDsMzH4gk8Y1sCOzSETMhyfwc5JX2hd4WU+ohyISa/Sd
IM1GLgDzq7QdljSmQJeWxo+RQO1zAqRBhFXo0TPswGRqz+tgRDwD5Go0VFV9CkNF
XPVv2erR4A/DgFQYdUoMHc228M1aiC5xXq9bc5AecTcnIWduIwuxOISNVpOXCw5F
/zEk4w+NVG9AloIWh6i2bECBFlSxV1F6fq5OvUE777ynA+gmfvoGyNcWe8YlRBrM
DA3V945WCBjI+gAN24t55AL9rErotJpc6ONNx41ulNcHDAe1iMmLa3PF6x9syiz/
jo/uP1NimM4KE2XAYi259f0utrj9EKyQSGkw+SlFL1JJzR5WlYOA04wQ/yKqd1Mq
QUvmugs15z+sz4O0xD6cfFBGGy110SCuvmFn+N8636TRuACM6VLn6o4RDvBIqJ8X
lFBeW2gyfqCxhb5wVEc2Wi9kq/oXgz3NFAzYPj1o0OxOECjZKSx9KKJ5TiUt1PPs
DTC5nIfAvitUY7ezFjgY4fZZ7ZmywRZ9hukbRmD7/GclE3z3hczK0kk4Z8+OQNGM
fwMMYLjBvRz8aTNSMFU2utXFdiMmNG3tUN17xUIYngZUMmcEZhQlD+16yD4Wak9y
fFeUikAVAbj2t37xv3f7rM1i1a97BfNr8uelh7ZVcH+1dCFxKquC8xXf1AI5NXQM
sXwPCh+fVUhwXC3EymfkwuPnq8ddL3lz4OkO2sTKq1dHcZSRshi/3Y1QR3DwGMsX
dqMmzAejVkM28hYMcYHjmx5guwMoe5diu2eNMWvQEZqf+07tTvb6z7M33/MUTbKo
O7ltphbEV0wf2dbJzkLC6lSP2y+EkaOYSSS/IyO/0u6kgjV3+5aHdZ4uxIJbTO0D
elRiRvxofMPDX0RQKXFpaYSkIlZ86/1unAwhfoSNAClk6AQPvADapnz3YBTTRivX
Vk9s0vvKynZqdBg2GWV4O9NAqWTbjlVw6fvM0zlkw2gpAMiXo9AUaTQfx9DR4Aco
XBipy8h9sAPTTH6gKSVoJRii6riafUo1+5HBqTjRhlvq63BjFQDntqmiDXrLyKPO
HkIFh8I+4Rgs4wboFMnRnH5FyclKTD2IOMFlaSLCsvKUEYFKxxLvlYZGUZEm4N9h
G/En7Kw7PiPx7cUC3SEGtcAyDLFrsCigYhc33kqeYJsubOPXgfxAvK1nhagEoeFT
HdmJPCsElxuwGcGsyzhgFvv8pgS/ZwcP6RgbbEnH58G0stfpA3iUt8LvudqawTzt
Rg8PF2j+ZPaZcoxU44/kuGBgtL2nTnlpLKWqCVwRtCySCmuZmgI1z8JuTG+M5eA7
pOFMjNaydrbA7dz8cfGiOjRVljtWWNHwSQbTtArhRHDuABm+IaDcDFAgLYPbfICd
vXfvemNuExJgEsgGBhdi9XegTfqv6SvGwRvPW5+k/f1CIrIMljNahZm/n9FE3TsO
ITKSuKSJ685R3p3HhaGTRZokKpsNXUr8bQ5/0HJPjoM6jxIrFJ0ncrV+/cCQywXS
ckCJxg3o+H3Axw73uD0l+L26G637jnbmhzyy06/n130i2Zvnjc3Ybv/jMCIYatH0
aE84odTnsJtETH0erNoUhpGmz/NMtY4Gt8L+MS5cZkIaj/pg1lWUK+qJAO1rzPhW
EmZdxx8lPTLLMFE2qbu/nhZC4NkO8rFFP8DvAavAgJ4PxlIcqIYaaVKJdvikx164
+ZQ9DAwZ8hY0yoyZ76A2kdx0wF+RudSGuDfgTQmggMAE8ZvzT+LHbER/4ChQdtZ9
cTs7I1IiA/ChrNUuukXFqUL9PteuBjXf+L9PSS26IenJmu73edd4fxf2JxM4eoZN
HZxHYR2c+fjIE9WpZEGK2XzbaNHdKJ4WHWkbXiHz2Uh77GyDDUY2uLbAIHE6i5lT
spQs9h1K3MpERj4wba0qJvuRlYS4wx5HIpFdWJL4ZiPqhXPMlNQozMCOyNsswo1l
bKhU/mPIDzLYggM0nAHIWSX4wj1mZ7j9Ycbag7gRALL/IzspBj6YxkhfmikJRc9h
vgCSNxYCFV7IVcv0BlgwwAyyzUxcUh8Nt3vyyW5/QybNiUP23uj/lZsPum24hqM4
MLXF/Dpw2FKusvwlBD6vfeO7TN47DTp25QeWQHAZh6veWSXKpJax3HH4ZQCvB2Gi
HaV3NjpG+s2oyaHVTbWTbu6i9sA+15vrn5kdM3a+UyOvRIDFW+FuitTLFwE2g/pZ
QbIhl2fMLTw3mp52MbIsJSzUZpOItqPANL68jD6OyN+6M2zuGGZC2aSZBCk06B0a
TgiUIbh13dl7a6Z91Z7k8/ke+UNgl08pEjCe/YWOB+hbt5iZTXhZJeiq9lLZupv/
omuHDAV3bxCPTALEQMxIpXm3b4aRO2ybmTpdT7BhkGEkkreDO3RxBjNsocFAz/im
Vg+/5xik+ULY2R/4hgyF6JEvTO+LCLbjWcb091yzxAH7chxUWNu3nnPGDefHmqCJ
9z+U+GMgH+AfTzEWkkbO1IYUlwUesRNLsd+JdcOzBZjbKwYUOGEGlPgNmCq0Phh/
0mT1Vz/ggpnETNceSyv1wC5Cb6U60Yxzz0C4SeOFWO90L40N2g28c7kd/JRq8ioV
xDa66MUod4zBG6QL1Tv6g6eni/2tEly3DHbPsxEEefAOFRc7xBaf2sBr0sgV0jF0
dRwcJQoAo4sFv/Et/2CosHL2JFhsRohXLk1w2GlliWzpx+hPTQCmWKptfhlbmV9O
SEAwV47OD379oykWhNAsftFb2syZqUoaCva62j0ILuCRf/15MS3vE7SJ5qtAcibi
kCIfCYF08DN3fp1U6+QfpKdyD9/+9WU4r3S5GfEaSeZWRWp53PDrWmmFUrbz7CKQ
N5WWfFhhqWbmqLtuif7/SHHTlorEdNdyVYDvcbT+feSA2aaizIZPWmZnFJEO45v8
5VXpCBkjnYJgPVaG/agkqM/lR3OvwQ+nGVL7A6ARU+ol5URGiO3uscTSU8LsTbXV
CAiDyL0z0tskLkbZiqqCbU1WAgdA8wZPZjQykeF5nnMyIG/hx+bdteCGpxuLTivi
VOV/DI23TBoukQSiYRzUO0of/edu1Yobo6Y0XGMWbDkcSQHV4cQkaVhVbKS6aqDP
sZga5ufAvaA2ffWxq+xg8efFuIv/gq4wo9R3eH/M0KIpWfTPI+zTK94HCIb1VbPD
eNYDhRGEVWfYRn1LhK0kIMkJ9bjfYTlFISzLLHbx3Q/wERlcSfHY9OXSLa7ssxUu
Cw5GXlXtQF1SnWIFMmjoXiCLnu0BtjrjtKQVu6+aFcfMHJkN0FbLR2ulQxSYPzJN
pP4qsckD/lZAczmgA0rruZlX5xbcVaXi1QHGbeFYyb0DlZMeq9e8L7ItCMl3VUx2
Xs10Unqd7tLkYVWkIgAmhSv1/FU/88lRqeXLbRbrOvDyZIuGYC8PoB/lVBTlmASg
CVunC5Q7JC1hyemwem4cqXd9lrszjgQ5RNbrXeCMiA9kJvvTw/psOIUvT4rrwwtk
I77DSSihY/L2VJbwZtMsahXFVpljGHpFoRsncDPMzydIcDGEvto/vTdIIfbr/65I
zjOvnVVH8WOqyRY4qGjzaLC49A0j+OCATZOP4R6goiGvs3kCW6xg8JK47Ctv+io7
q3rCagh/PuemzjSyNjCZLUh1E493E1jaoW6sUe+I6EQNn1MHPC2h5GgAy/2OrOQk
GRoxxla4m9a38ONrnHnpaRxGUMtM0JJTXfJ0xlk1/4ciRe9PbcRhwPpCA/K7Yho1
MgBMr66HypEHayV6UcTe9B3ZsURWIM0G8kNhzzH73R8l/MnxDNJxiiCp186zwpKu
WDbbEsn+vdeNa/ioLb8Dn8qzCr683AJMwGz9RfFJqzVBeD+YYCgIC0yHuFcT5tcK
zQ0aqtYQqDo/Qg6/GpHycsp7S31ostZDIdj6IfG+71HQBWgXWKDJP1rAWAFiCG7M
IUdpPbtw5eRYRZGbWY5yIFOoTKuIOyxj44w+s/4YTiHxrtEcwPCJglLMdIGD3Q9h
YZP9WTcteUFnTf76C5InVkav0a536/kDPTTlsnvNkOFk4vsW92X9Pqaia0BPNCY+
HOw+y9M74ENhCz01575D8JqvQyrOMTfK+E/6qK4YdvZhksdx1janDFr/CbDlBHEj
tKyaTXlTBH8ok7CE7DOJLH9d3Nws1DkQJZ2ud43JCX3CCS+Na5bxyJqx9QeO7MUM
lk/ePzzTRePjqwBsUziHioH0OywCTzOs0mAZqGDEYEsWlK5tFGeoU9waU7nQ09Dd
34V7df7fOplkUSRfmALDmZERX9E86Rnuy04ZZoeClsPsEPze2wGnLIMZD2I+DX4v
C9e78OU+dzEsdkmzHcoAk1UxVT3FmWVPPBdqMqAPCKK2ji82siQ7B8obDu642ZGr
fXrcTg54Lh0CBLeL4O9xbfj2lWaY8JNBjTZdIGB95+DSeyDwp/W1Sy9i2rPy4IOF
esmRMZ1ZerMc4d0fOuZtgjqCH7/3+sBhkwoxDDJC0wltZlg0ls6Imj+C8R3Oz4Ik
ccDvKnSqnymaL+VCAQVv4bwrG+Jj+ZUzO4QtLG5TFVpLw8kS4GCoB5Xi7e79gwpx
fdRW8mVFX31T2Q/FMTZlfMyoajDTwpzxjffqW4RQHE0j9LaZmgMG8fVLE5ZikpF4
DbWUfaZ1vCsogb2xqGoZTxc8gllS/EQltyQx5iUD5GOC3XgvoG3bEMPShzgwsw6r
j8KpLWpSV3Mg2gbRCS6Y7CbaTX9YU/qB+VZf6wnAHcYrj7QB0/UM7T6HHfl6bWQD
4vdPOAHJuLKnbjgneLW6OMl/vv6UAh1xsbFYa8mgw1g9KmzX9rPMoF4Tq675sGdU
Wb2YsErIwk1FQaBI2yhi6qmnPEUU1HCWavomrfN1ugzcEEqu5AQvBFUlDHugdli4
YX204EJEuHO1zuMAnAZ+wF18mUh0AM6y6rVFHQjIsCRXCZPuC7YDzFHGIgKwJ8as
jyJ+ropHly5YXdWQq8/pmscMSdr/6CZXdeE451QVBZzBD8pPJFcMMoY+dirDPujg
xdXMbJpeirF+OEmPiyR1fy4QWOr4EaZl1Vjwa1v798lQw4vBKhp89E9Bt1VMe/EU
gBJu7pmornEEuSa9y6qi8c0UPXEHZQ9KfflCDKA/ZnDBBK3KVbbCbKGaCqey0vRO
JS/LWa09khwB7Yr6bl0djUs9k+8TvIyNJZylx9utryGOCSS4IGU7YWBEMKw4PsSd
KvHqTCM9fPyPtpC2U99VzyqSPY+CFjrGl9LsBNYlQSbm1PD0z87+hHamBDsUbTh8
zrM1Eikx2uhSyz7lbIelwW8zbZgf5s+9Oy98TB+1mAWBdGBDzUGNgOPDBC2g2IHd
5/OiSpvRyP/4GnI/J2TIrXeAv9+eu+TMKPWejz00FpjHf899WeWSIn2rGK6oo59l
uBxEvov2jJE3/AQLvzIztYNsyfedO8GVqAGmzgSLgKMnEkXpk3yqCQ9+gKfPnUkJ
+tjMGvHRSmQSxOPL1iEE5Ccb88eMXEeYOIMN85aXxeLSe8YhxIBtM6qmSPG6Qr2O
Xw/sybF54GYgvfnQh/BiDB+up2Ob9A90bBoUvwJaIHjtvqTDjAAPEFyadWc92fxq
+YrsqGr5m1bN3FZPz44GDibbrohpln8FruVKILfubjIdjgLnF/cEZ397ExRxldvX
PPlVKdpYUjobrjKNzstuvsrIkboO8hOi1w4BjtlgL7DuFQHY2r9G+fLa82+t46ZN
bKiRzNm4ArW+OLN5AEYm8UGEc+dbY5+fWtpOO3d6P5Tijy3/VqucRqvesELo9R77
fvfN/CffyrRCOD8mFp9Z3CNg2zm7RREBiHaXQLKt8hBD7iX/OIavPIzharsnFz+J
6UhJQMtV7Qc1KpI0MuP4N+8h0yBhuIPMGlcdYiGAFYguWtmsoMI/sCfeU6gj1C/g
iGAKFZs6tp2ZvckC/LLnZ0lLv/rfxCQag+OH4TW5SLOHwtZPk94k/NtRDCV6eH04
0GlguVN1csGdyFT3nXimDTE5rIQIzZPZB79sliG631vKntizbv4gXmefhlmWkI2L
9BzH/l8kon5M2gLB6Affbj283/kKXRYXvoIAMHSd0VrBhdesXnlZXwKmG0ODU5Pe
1zXoTyQAL1tx0Eyy/xGmtgKJfQzFfoKynCiii/a1FZ3e8gyGjArDi1/H/vXXZQh/
ZzzxNudqN3Z7kCdH+UfzMiCY0zFfVw0NGDEk4Rx/lB1lQguFv7BYvrtt2dyxo8Mx
J1lewdj3G6wHj3NWADysH5ipYWy8Bn2Y3U42/MUXhqpijjWuK2TO3qTROZUHWjMr
Zhz3Pkwj/V+Csp4veat25b971nmtC/Q1pjWhMIl3hN/8Dysh80JLYS6IxTiq/7Lq
7cOFWtMNSPSe/yod01uW80qeP7spemZ+FNGAh67qykYTIE9ROBr67tbXcXc7IDMP
y1aA2gnc6nT7qdgH5SwK2nm7iFk+QN/Lvrzhcx+rh5t5kZBtHe84DHWSKUQTgmFl
OmNggcNdNOA64zwtz4VlO5ZzTFQqCLyL9yhdy6dgU84VzVIY6JkA/7QO+SL+C5g1
pxNSGeEQQMP7rO9MBpIKF0m1XgjOxrfMKxrvBtDabAs9BHpTsI9xBxdqjwfnK+tR
Dr36+fk0LTcG0nLzGGqygFtdpTbTZBN7JtWD90SQFGxQ5xNPwOpc6tUVQIGANpoz
Te/lqE3e9m8s7LqbCHqfLhLKLbmyDVJkPYsFj+9PvcOgwp+dsD8tYt1sPUaM+8nt
04Ec6d7dD4AzSUfUTsksRzZIL8NcOjzcj08l1tN8V+onbvwUZNzLnheMtK/zSabv
luxex0vm5ydnR4//6crhZ6vKNSJbhtQNEFIrBG6RM7IM/2v1+YVcIdzHogc8cIOJ
s0xYX9qDqI+FZgdwgdbV+cCHUM2Nglu6YVzYyoWOH2dEm50XT25JRkmNqnomQaxl
QY+vA9xrqja48g6j1ZFgNrwJt1UeAsxqQLYEdD96siQFIOPEwh6K0KDUC3B1AgAM
c2pWWgCmLqBJoWzXabRyO4Iq5Pgj3igWkPwoe+zKvW3FYKNaWO/2NPtzIl5077P3
75o+heLSJzpFDMe0o73WSo60sUET69Dt8gySjGx+NRPb5jQSebBe6chycpay/Tur
r/auVy8tJNzNkvvtuuw92/F3Gm3/n1y50q+sUE36YdhfMXy5ml5vkU3cDm92znSp
duNZaOk2xmXMK7qcBmNsxyQXY9L48Pr+drHR8GUjcJFfJHN+d92YZO+E2sOpF3HQ
VAhAv1W2oKf5rXNuwPS2EJ+97GahCcog+9ocLJS6U8QJi0SRuOTNhZc4xd1b4omE
RUZQGXgSJhYYt/PUoRPoHHxVc5lz0xrHCjCLokmTKjxc50Q8VSfKgZOpRHgIy0wT
gbPoVTmU1jTHtU73Wq7oVfCTPl/g4jXwGSU4w8p6Oqdkb41TXVayAvmb4Knbp0iq
oUtI7nG5A57PfYajs77+s1a+V5FVPY9EnE9GCBKjZfIHZrDFAB6crZcSdz28w2eZ
T94PCcjM7S6fR/uDiiaTccgipkRPDtBjcUY4a8bf9aV1PaSxwiX898gaH++Zs5Km
kAsB5GZ0euc506j0F/3EDez/na6hDH+BGVgb4/NnycI3TgMRman4/TNkdrKJ0lag
lghNdbDBsvF4w/f5v3f+aqCtWQk2HUNHR8CyziLYVkCKGWyBa4gXDncoosLdMqwk
4IZevkIGYlSAIPs3xtgolbods8TWbGr/uGrO0r/ahwBOAnoHHR6RUL+guLyAUZXF
L8zeri0nNQIp9gciRDZ6Q3Oe/E5PnSTDKLNfQHdFOO9WXzdWmfQnZSH6jo5WlTwQ
s1ma0wUFtKBrejdKVBC3oBZ6r08dC3Bnor/1Cv1o6nly8i+6l8c1zMkPWoBGKWjE
u8etYN2XljUqe6qbsV/MTN3l7r4aleTLwcSL4evB0mFcriAwqWQ656H9BzNLjQbO
6Tz4zQ37vNi5WA9awOvnNuGU2t6V+jDeUQn/YN7SaIlLezTmvz+l+qMhRri6e/mi
oXpAfxbPuau1CEx524fy/XUL8nl9RJHMf+IDd3fYzfXVR4n96dRRK4sbyU7ub9cc
4ImtpnWCVBw70/48JBASRReHu4T/nVtIIjSco1zQeqCZCLC0kVcz0/oI3lk2tfdj
kvL5QTJbd2htr26ivdJLR11NuOX2zIi6XyYCXjodTpYhLsM+l6Mtj1cLes4wDEiH
E1jmAwVIgZtOMJjgYmMY3o7QVndeptdowq11ds3xK47H4H8J1zdWBg5xlIJk1LgV
tnHqkyTI5qsX10tmNILHf4jk0Pnj6OCkQZOmLYa/ibvaL9OWVuaCGb6P+J/Vw5Vs
wTv9BQ9IY3KhlmzRziiskHJVHmAi5K+UD4fnDyyfCFPGIaVdxnPPUMhywcsCy2JP
G2XFjAdR/ZiIGssnqCXniohxswhfX32kRVHmvMaS3ScAsUQk4fDec6EHJzOlsnU+
77zp7g4ITZHy/nikgx6vbtOxODTTdRwmiI5flD0vluiGA/urSUCxwQ20mK30dcKG
JRsFx6dgVT5CPt0OaRS3CwaCEOb4EEZlkaCgZ1FmORsKHGaw56R6o0jVdClVwEEN
xhdVpoMv1H7hyqZCn7C+A5KjNMvW5F+tEzdsVZ+iBq0EiydtFMzrd2K3AFnn/eoP
bB8M5QJ6MO3MZr+OWBNkL7+AcjN3uRLJY99a+tlBzEqVCTplSUjexWN2N9ZSgp1I
xRAWRkh1AnAwEEgN+G9/RoRsby82F8VAKD8SjFOVh2gtbU6WUl10r8YzIEkduNiy
+EBMR5n4uYQQNgHEbPz8V11GNHavMi+B7ulOmo3aL4FwfsM1xlsnwbC454NGn75Q
duDINk92GpH1Z1CDSspy3QUYjcoOhOaHJYf2PM/NICYO1t/2G6vu5jrlT2CKdHpw
FupcAYZFNQfRG80/PU4wYM6eVLw4+9El3TYFWFDIJECE5emorQhI1TFR8d1X1dIY
9/x5r2/ArOWeWwnoHZgtU5wEhB+1i6nUSXpMp2KlMJzjAeslJ24s8Uhpp5g1q+IJ
uJBqmxNrXmILRFWGmj/ohOQzT5EAv3ue4999htx6rC1lEz164B66D7g9MaPV6Z2H
6yjiVQEdrQzHOc/cFj7sKzgauwB7r2KhvIEe2g0vpcEXp6PXQ5gqE5JbonAI31Q/
XhEtmslO3CCOKedGfVwcsH69NUqznsxOi5k7cAwxwg7UR+VkxIpv/PnyW/CERiFm
CYgqG4rIxnqfhXUUMwXcFeqslPAqKgsXeEzQQyEGJ1WaBKOAvECw4WbnWfgDtIRR
f6SaQMPJUCm/ebos0Cg0x9GkqQEs9dn9aF0Ugvu/tOMSKALClhiCmNVjXKlBizvt
kAFIT1M0A2MYonXkTXniP0vc3OGyuRv4XbsMMjrQbgqWjFt+kubzEtIgSQ+WhVte
Uno0ShMxjwIqOyz+WXM11OOt4CETF5is4bwhVHgiM0xHwcMBhHlZNdSTgC/kddy+
T+bbpWAlqdQgo8Lxw4nfPpSPJhQk4TTZQ6nWCLkIdm4ghNFZEwR6bQeXCqHPoZY4
9Issq64EkzFFNH+Xk0B8e2mEWHfnoPv5WzifRVTfn5RxedXewvKPGsf7l/DQlpYr
8fwFJ78S9Rk5HgYOKmjMuPzXQ+Y2ElvNMzyVpIFAVlZskOC+QT6526PX94cWZuK3
/Szn81IXstdMNT24Bi6hwMS5xezYQfC5s/JQXEyyzDVohf+aRkXWh0n0ruP16vLY
hCHyhyRLc3gR46sOOvXw9YmQlp1ccmwhesvu/mTjkPYyCZVVUD6II8r8ktiL2JWi
65oFAgmVaCLb2Wf89DDJgMfcXZTbBAiwtJ1n3ceGTQNOvvs/cNEWKI5h+J5cMEbI
YAlmKZfnmiGlYM8XMoQdgfAUwWtLnvP4N3SnxMiANsvAoizWYRXaSy3Zjf0Qm+V6
Y5zOvSL3cnFiNBwaYhmuA5JBGAn4HcNTCBNlVo4jAgEYVbIEaEq89Xhk/DpS6R3l
P18bIP1Zmd63txQcDFZUqkChaIs/G1ZicsblSnl2HqBUclNmuyxxN6eGrwLSEDs+
wGoJxVHEm87ySTUXQluVAE+gv5lB0QsSqpqc7qNx0bXCdfLdNs87a7oQNvAdRsUr
QV3KczkAXWpji6DPMK/66Vf8c9sq3V2bDrJEZcKHxG7Cr/5nE3aGvr7iajAWvEFT
rFmtSKeFBdQpYdA1E0WlQSqsHIG2AyN6X3FS4WwdlQOAVubKqfwnANn9WNvkumOH
ASPqyhy0r9Z73cxTf/mlhkG67MOfRxNHvyeSK3lX2+NQT8I+pYTD8AquCtf69xnz
cLkn8gAjWohx2htK5Iv8Tf66QdvdPqxuv6TgemkW4T+AY8DRTp7zGPLN0j1qq1kA
6NVnUkc4STbKFc/toT0fZOgkxZnA77SsPzHJo4Q0xsT5aC9uQIoPok76NvN0bEs+
bUkiFJw4aJd6y/Mvtv5op4S66G2Bi1tzuuiIWCkzFkYYLb/izc1Yr1n3iP+mgayo
QOCmraCyXGJRKD4ve+Lw46Mvd5OQAywnPMLfXVdnUtVMtHUFSC5EfiWRxpMQBlrg
3ezBxABkteLjaM2J9EfNcL+1w3FRZSLilP/Zj/FAZ6e4em1mjYNEekYSRUXLqL/q
3c5ji/EwwFiFpJQYP+uZ9CTdVYJh7ILN1q+9qF2VKJJOrXeZ+duRQ1N5tUcUuhRt
UOqEJgS2aPu+/sp9zoI5YTvQWindpgc8O8BpAtYnzm8ez92sHTUB1SEeKWqT7tCl
vkqarNhyDdSjK7xDGFeRDueAHZbIg47QkWbZQzEv2F1k2KrhTJButMc1+7LyAExs
NrbWzvC0s/si/SakXoICJ4I+m9qvamQJQq7MNl/CxxA3oUr8AYFRoyP3lEw5VT5p
EmoMFbfJFQH5t2NogE3n4dSwpQq86xc5NEi7+qtOMR3OXcyfDyaWddkG6Tm9VGfR
wlxhm8F8nYtKSWryZMQOsWz5wyLtxyS/E5cJgXceDNWY+r/cA9JGTcHOjsLrZXgI
0nkuLucqA17ln1BSYjeAitqiYUjQTJEl75rqFYKvBRpEz1qCx1ee8HnS6NgSXtpk
mnwrMGFtg2YfsLREHAt98sHyVBg11yv3384NLpk1SG4f2XRStzzm4cP4JWpm0U/1
Qs5R6madbocmF1T7NHH+vJImquMx/vzBIBIhak1iQzJ80zOaDfAt5abNtyTOeY51
2p9P3f/vbdlKL2REvwOh5g9kfSe7hhQIIs5CLrXixaXwwHELk/XAe/Fz+klyhKhv
UtISrBYcZtf+Kp8FnKR6f2iUHYefOAvIoeA8AE1qODhtDzrLaH6ZBK7Gxvm+guYw
MV6FrOiJCZhuR5u85VLtuIpKDaQCLyP50grNsbFKvWvwXOVYdvnximYgWxur+khl
n+Bavq5Aete6qXgT67dYtmNUmrtvcs7UQUOHddcR8NCxjqmJBv+TB4+evRvVWwbi
ZFmW+9AHlUg6i5WD0uX5ieoE+1Ez1o0GWsl0UA4JziCRXBMyf6hFsg9YmLa22BNK
7VMIcNIS5raXg/SLxVHcN3oipqAIu/eWK7+H7kuqGquD57DuPIS7TsUk8XPwU5Oy
F0X1ErgSJTicZP5JYnTI3UF+H6s6mCXDO1HKGV+yqcXfcaqecBr+07WGd7WGFhWs
QG0md/hB9YcLC83bE0OQAuomD3kidLvV3hy9XVgv6sxkQLQuLusloaSDIdCPvsVd
mQiuQYgHGBfy7D/On86vNzyRpQCpvIqtgH2JWuW0J0FGvX+00YSFDzlutM7z5CrE
vLfs7bCJ6FYyDowCtYdCYrTa9w8asW0F/33XEhMllRe0vpjaY5hzna5FE5wVQic5
rKjxQHmw6eQXKmJ6RE6QvtM8ytg0ilnBg1Z2UUuuwHal9aOq39wRktOXYeXx5mWI
dBMl9T33CDvqNWMdcePYqusxt4ZIj3U5HESwzAE8FxOZN28EvTxfcUT5GsjqXRYQ
0yOYlNcI0D9W7K+aaLcv43dujlaO7CChv5QYN348XLKfhiof3miAkyeFfserlMWI
NrAVptxkSjpST1GAR923UGFK/qcLzU2akDJSsGI9w7He3cwYMtwaw2wtRPwh5PAc
SP7OHYTALGsPUpN5JLshlR5d2+AwjQRNXgo+I7kn9sSNc52hmgfQpRvXc9vRYBzx
p1+6ZU6S2TFBzLJYbsfiwKZCikYAi43AfSHIC3Im0xzqtAhVLqea1tz2kMvmAc5n
xVrIRW1ugoj/FpVDFunlf7H7Ldp2hOGrG2bMXrOcQ+byeBpmKliEFvs+4zYeWYuk
S0XXY0Q++tyMThcCxjHaKNvxWRjBkv5LhPr8CgIGeEYcZpEJwoIHbNWDP7HY79fv
/xl1QOZKC1z/DeJm7zN/vghEFJgkTmbUP0nQqmADpGJEkwsb3ZnKK+1/34iw/A85
OewyVB7VONqQArBz3MhaGsOd2C5G66GaW6qeV4l+w7WKFS/r5hBcBRE/L0lrqu5K
jFJZ+/7nSg4WdPtr78Ves8JTB6VTNU0Lt4MlaBWdxdHoWuvZRaWDIH/OhEnlp+YK
mQcjtZYwOrpHIAqsgIE6IUhJljfpDu6hgZOq5hsp/Lhooq4wc3I/SG3y9Dc/BlYw
kYLOm4QIGZDztC02uvBshHMPN+I1htpCqZx9VhPy4LE7I+ovW/mKnk5kh5PxVXFg
qsUl/y+08hmG8EWxME9J8uak+bSoznBSamdd0gucWaphb2eXgUSVNxasHcHGebxA
z1IhFlrfpPsTc14CXMiZENY1pFwYBCtLdkhm9qDz/jNwi452SMTotUVVvSmvyS+b
1BhiBO6uIatG5RoFc3gg/jQzPiGrtUX0EqLpHNYCMFUhfRDt0ug/AJmSPqnPNUxK
lY1E8AtZ6qWdJV2XC5fZkDK5jyNEvtjsBaJhPs2a9vGHJWZjQJnVALyyswAxBPzO
usdIE9W6GKNMUKoZqbsxBZdQyIc6mUVOmPCV+mak0RTgP5GVBHj/8R3mv+sYiwQ2
IuznKuAWu7Xzy0JzkXHDasy5IbdC/8N5J2cSKEzwnmy+JDR7wyH7oKefOk9dDyUR
CHorlLmN56drAt6r0sUugyWbhzveU41lsKnko7gYiD0SZktxMmslJrDq825d77xT
yBv9TJzg3KGK3iRx3dcX3I1wHYlyxytrG18h9S7jJ9arCN0hi2ofOR04xRUv2dWQ
dfn0IJ5KDDu84LrlWcj1J7+ChDv13YWet3HNLHx9PxmltFIMz0RPb/zPbTt7To4r
XCRTEcd1PVFttvv4oVv1XjYKcPUyaUYZsjH/rnCT5L32A9Dbu2iujCEDJP44iRI0
haf2WqBFB/vZ8URHgkUPz+dtTH5P9ejT+a+opGorsWYSXol4fSqhdIXezELcla1t
Mk7NXLH67knx3vPmHJu4MoqQGEDnZgROucLxhA7488T5ozKohw8jgzIvAsupHns9
hnrPOcVXdTdAGAfaoWh5HRudaAru+7uqX4WiEj7ZlV6dtfyz368XA6Ha0ipO+MCh
4KB2M2rCloHqDVoHkrtLhwYFuqABlnFJ3o71brdl7vA1dCguC2pzQn+9YIi9u2ql
tIrk/r8hyZvsjO8vBgMebFhjfaCfERT72HO5rwieKG36xlz9UZY+52VpdAtbnTLB
hEi9JBtK6fK0txRYefKNyz+JPaehaOZX83xjYuglyXyr2yDUZX6t7tYdLMV+tG13
maQS/xkZS3UGaLFwIh8x1Wr307sGqfGKsvIuLnL1tNhavhJipbeQ4L2/d66UrbJF
uSbCPwRV7yXAnE/rFDTLYXnOWXWrWBDDwsjfZv3E3k2q0OOwQotDLj5PNot7KqQH
r23+QAGu3H+Zj8tSd9BWXnAZYM3Sjcb6inch5aHLdsWfZTD4U72MN4PNAwNbOGIy
x5aHBD5JPUMXKo+n8wbTdQqoiBQsEN34B/VxyPX89xNnLLyl26b6wRUtZ+K5u/jK
wtQ7FmE90wWzgB+UQ80gDc0NB+nHM9RmwiGbOZXdoVabusnnaEckH+6F+G3DYUOh
F3weaoJCSXFSyFc25cW6J0bOVLXwk8KnfmAYfsJZVe5tuUmHU7GgsuvuD6Jg/c7L
1HiqtfICQQPWDw9VgiuBfm5irIJABs6OfqtTgiW7FEpkMfrmHSWT4SR/IiKDUjFZ
dcCt/6JWZK2kHgikR0A2RykTyYl75LocLlMxCDOdZcIhpqELgFndoZw6mvR3wWcE
/CMOAS/LrDRPCOCmiDOP6LX5OrgHcIwcOu3f5a70pSReWpawsSsA41wwzbsiiHEr
qkQv2WaGTEu5F3XrkhArWNvaQfniljIwMW/zeszh5aDikF26RlN2c6Aok6wGemMi
Qa5P/Dx9w+77WpG29XGFmq1LyOsRa5CQiyI163zhn8hia3DaoTmlEJoLMG1G132Q
h0fZbuV5A+8W7Iz43ypvZufkiPYSuxHn4dgAKqFKbhFJDFFvn4QAmYB0HVGPrNzM
vUpHIY39FtbTYH38+5WXj90Idg85+ab/8U7vrCzb6TCQ4XWdXtoc+u1BU99s56aU
vVhQwcxnDcYGszEg5BbJkBTBvmjKXnFtOJcDERIFQomguY3KC+EsFF5r2UZCVPT2
e+RFh8k5uO9tQApeig8BMRZzJQyF1Pbr+ImIwbWAHZxcRj/ly3w8/cS+M8y8DxVc
AnmQwlDYPmaGk/fwDQuYDX7PtB5XvRqXSDJ0gtjJqGSByNSg2QV5B//Yihnutg7M
RBJ1hi8/zdJ5gz7j4nPl/gGMT53CQRNy0lDdtT6qZgdjAMQrEprrdUDD7pycYG3/
KJVEvZyu4RcuYsfpVRnvTfH9SiEZQJhfReUdm5Bs2a9M/oLC5qTMg6OF0RDFnVCL
8HNkyXwx5yLsUycomiRkyZX6ZFrIkh5dsWf/kJ1XxgnbhaoA+ojXsBe//VVB969D
Wdv3x6UI7iUQCN1ZLywsyQdt8mU2BzcEqohxYamJnwTKytbSHYExmVMBgwVcF0sM
AukboHxbHHtZuRamY2324etLwICMj9e4WH5tGecnLQpMaflLeG8tE4gi2B/4dLDo
8ogW9pRH2CCQktOlGhB9KuFEdK6+yn+HGiSi216wv07zrGwHjmXeRL3pigh9ZzA9
z0ZP2qHqGUzGRx+NAYdbGEeCgXIA8IOmwZrI/n8Q2mWw6BTwnG3RjqZV2QuCZkSg
EM0Tb82ps9V7hjISHjzZJkZsHqS3DtJwTlRqIk7jMYIg16CmiMYD6NPVQ4xBtuL8
1EAUVd2eN+cFUqqCD9koqo9hZWkox965sEfjGAfXx1DyvgPz1//cVnUjGG3zzHNw
rlz2DkFfFF86vkQPjUP+LGdZ5HL2VTP+34kmTZP5YNgWHxWyYE2KY/XN86bv4Y7o
h9pN/rBg51iSyUBPXVmnjqQpyM7uwDd54UpoAYMOlraV5G2VzECttva4JUibuQW/
+hcdkAaev+oCkyktQGAT3UK+MYO/dhpt1WY1Dt5S5ke8Ejmky8S9CZ9W0rXHnrbc
5Hit5a3MADkzcuqTxpiw0xC8RpDp7iColg3yJ8vQpe5OPgyeDrcNslu9QDldXNNE
RXcKvBYcN2fjQ39UvB2RGFqbo6+cq55TqXfK1hh/saTVkApDNog1oyR0etXXnA9s
+xIDq6hhx+w1s3c6Vy9DkDALjo93ASLmpqtLfZ3qb8MK0TAzcqsYyzMang3LHn/S
oa2PU2TEO8nlTYfWyp9eeapYMcc8HUr5XbudNpxMXEbLfuigrF8MWi4ljz8elbKH
QkJ2om+GT40UP1/zGmVLfXsQ61IqDtVZCtlzJhuGsKZ/3xJfgtfAc7X/yx9yZowX
q6/Bjpd9VJClLezxYQ+g6w6HjdUNJ06rrYke3rF/FfF7prPlyRbsmkAt3u8VVYrR
1t3yGDYobnnRKfL1NAiyXjb0T/iVqeiOrBPmVE82b/iEd7yIIm848WJ/ur3ecD9y
BHLmsXZ9/fa11U3pRlNUOJpNgaDTjDrMEFMvAe7pz06vaiZ0d1uaIbLFO8/22TWy
+8EbParQL7Km8MbUupZPiBFAlG1K+uc6RJiZFsK/U21xrA5jVdHwRdf7lApoXlgk
ApMWzNfcwSySPaToBTFNVz7WuTgDlEp4gXX8yVN0YwROlvj6Crdhmh+WlUgWVjfR
a3ppucyj08ooQ6tAoblBArR+RMcBNz6qArQMS7njNDu75i19vxqa+RwMGwnNlAo0
Q5ydSoJHuZFUEVd33c542LeLGEZp4BN68fZHXwArzfYgG4O0hmb9QGK0xt4TVvCx
XUnm0CiQZd49jO3gqmSLu0fiLnOSeLUIvUYc5GqDIU/v8y3fozrDAPN30WJZzC78
foLjZq96CrLVKecf2fLUXp5+CtTgz9UPbqPfUAyCHhWGhPJbK3THzbodHgjHd3FS
Gew+AB5YGct9V0ml1kZHo17AapKa6U0DQFoZy7lLYnuhZZG3dGifQR43DcK+RhYg
8Ou1jaLXKt7UiPj7ekI9wmkotP6yuwmSI4WBfpWXgE3UgpReCV9PxFIOsZXG1Sa7
l8Sk+hV2TmTfQPneZ0hlNnTgjQF21gzxnxFoZTj6GmiMXSv0H/OoU2R4vWRMwQBp
CTGi1lixolQWFl0M+1VCFQkLO1l1bGGNKecyV9x6hIHqIpS0ANo8hJoc0EgxQIH8
29PbTixikRX1+o/rye5nUqtxl9cHw9oGM3xaX+icFY1oyOe6CQFCMQKwOkGhtH3e
RLbPjztHDQgYg6z7/KYOwICLp7nwJHo12CA/jb+AojZzIzxH28nRDH3uBjw4Z7pg
z/AGlVzNn1iwE9TxHgog4dF7e1n87NnjPtCPPlhbBQ+TDcfKoS/YfdC1r6Qpn+Sq
B/tQOHWiJqow1WbkeFNALDrY7wEpYlguq90oTuGAwHrbM1EHFPG8HjPBBQ967emS
LYZTZjzT/fWP43pzO9/vUxjQsxAmRUUu3FA6S7C2O/hL64Znb2SPIAm+opd0umBh
tUxV0m3HyS+5GSRRC2E4Uq+7di0d1XLJ3a2dqRfrfCnidmlDj5EtJPedfyPiRLyS
JWnAqX8JaZwo94hIfMUp8sXKhKtmQD7aViENsofTIQv0iw+FVUa+dDboyAOk6jX3
WK1F93Iz6xRiCozAJtMX5ZdSoNNgX7AJ5YSc/F7Hu6qfiKoicJm7ZJea1zjXd/Ga
4ZvJLk9sD8NmYfzylCOTgZtLhmgfxSyKkHHewEjxKmXBAJOXRaxxvJ/nrxw/hICU
Atv+FKGZUnYpHv1ji/qmJMdTJWyGKp7YLbTqWdzONzrQQCCZxYtJ0YjH5lFMEB9D
wNOoKOjquCryD48lMi25Z5HQ9JfdRIJ1cfISlqq2z+m+yttjPK7pf8LVySAvq1do
DamwYHAjwis23WLUp0FPDBYgXPNJT95FrAM/X0dzZys78qxn1bno1X+0c27HDwWc
BwX65/BE5P7eDC7i+Q2FIxRzag3klZPVJo+MhJgUv7Q3NelrHNJqEg1fQMpJxqEI
4glWsEFUP+dRSVKbeMUXBn+MTw4tJ3dPtpAyKJ38q9bzNrUEZGm/Bjnfe/E6sOhu
3hHbmI1gP3U2eyHqYJAJ4BMSmGXhGV33e9+ld8P/Smy5fIPxSEAlSjX1fQQR+Ra/
u1RwozAlpPqRpjNNJ09BOjiRzqH8sNtpvC1xAVcwYmztzoRLZFA2jPmGt7wIfSD/
9Zxp8x/t0af7FVzkbP7HrQhjUiqJH28jaKuJuVhUE9xjdS+DlXpCDeP/QqUcuJXR
RlDBwvPembNPnl3G4CndwMFohgqxW8uvPxkdtFZiQsvqozpi8kV1t49xpCpPhXmh
JLHalRqCGjAUqVdeLb10cnuB6RSl78ay6Qk7jK0rSMAqrj1+XheR1w+EGsRKtuPS
f+i6e8vvxAT+X6RQiXMwTPiL8+kypiaz/dnHHxoJ2oezYEPpoA12rc7cawwOUohU
AiNdvl7SM/s8gE46QN55cx2ivw2+rc0qZG5bXQGFsLbTrHKcNq9/bnNl3e9jQ8lk
K1iS7be4ZRahhrXlWdL1SLOfGYQa2H0c1paEQ8+rJogIdiRBUB7ICIwdPvI5mTUG
o1Z29eBClptQt7WBRg5d6gbM2zihwpoAugEp3ktFaLu2jNXlkBy2H+eUfB2cAls+
rJjHf0ThQNekthQXlu8EDE+GON8Kh0M0xd05rsRZcMDLhryQpJx+OqkjwEKyFGQB
/Y65ZKypeHQMWKvdosTLpkfjnDbBoHQWqjAnmWyTr5mlvl7F4GgbAPzNOpUZ72sF
xpM7SAskH62u2OWJBkOnsgNR9u+T86ER/IdnyTh9bN7eyVCMMhtV7nBprATy8Lww
zP88UXy4Y4/JZfL7pKyX1FcgXbHsjGrfIa2oXsLw/rqNoZBg5zWMJd4EeTpMbcDp
2ADtRKvalNFtA62oKmhk0KOXX16uSyEf6SEHYNHoqDcVXueva124xXpYTsv9JTx1
eNs+SSUOcqCgCulNkppgbQUrYfpkvBX+Li01oRg6aPjYoaaU5xp7qb7/Mcua4VYh
HbuDfUwxdFrlwlhxvPCreF957DWLvDCb5Xllsu5LJwj4HSVB9VkDjWAB2kYCxlx2
DePtz/64/so4VF3/MsLYVeKrPVUmVyYhexyQ9qbRh2QcG3WCtU7rxNN7DbMW7hhz
lDArbKnzoBfCVoTxI3tnZsRWPkDMrJ/Ht2WsmiaYLjh5nL8wzyrl5aDxX23r5va2
zspntlVna1Oejjh4Q6InXe57/E9VIsuj+9f13wVS4Rj1+C1SUb66CaY5O6z4hIOX
WFhEqTOgYIwuoVceZPZ7mEpNF0kGcvXAIg+7ycqvkYjvKo6bThxKGtNiVP0i01Dc
cZfz5eEb6sb+r9KqzzN8mGbt5fHAKj+GIhSaSCXvH62lxtMcs9pRUX5s9p2Jv1gq
LHo9dMHnzprO/VVRE3OkbNYOxi/RkWQKHpiq8Xh0Tu1jA3a6rxvy4JVWtUYEEL3b
fva4UJKvijIUGk8BlHd4YDFPxlE7ecNb9oxr7b06Hsl6yyx3eZbinpfy92V3vUf3
qyLbQb/936f536g3fd1Fc2KSLRLXhHWRwSBi4ewHVYbpy3zHavekYrhczi4Mpu0W
0raa6kFRwJXJGr14jYR07Zg78jvxyVr0bCRM6akx6zdPHnFrYKWJydmc3OCQf2ZV
6uGlCK1gS/VtcMxhDRdDwfChBMOqFr6t+iWF45IO0iXrQjYFBsOKMBxVAbKzDkMJ
RJv1bAaIbG+U52vTjpEQOqnBnlUTIdxTQfytPP6s86xTWH/jERUY2VaHdhGvgK1/
qV4JGO9v9MrMXmp+DaZe6MDF2IiKmzKtYVHZRYn5rLFH+DEIChgIoIN6lrRXaHJj
cropACzW82ixuFgrf9TjHWOOS0Y53hLy4gSNiTyh/tkCSf6QUygbfmFNP5T1dWpw
oUSURco/jBWCP90OnfWZCPVmrJ5CcWpZnmH3ZOYWTKJtSzEAy1U1udkuaxDEoeWO
P/g2/mctxYazwjCbR5Z20y/8QeWoP9xv/iekCJY4pBR730k7lfiu3W4JQusEVAui
XKqbwSYnhUt9qhBpxCIxM6Ny18SPXsembcchQXAk7Cm7jNtTA7gKi8sRMcoJC9CY
Y3yRuFiUtb4Mz4TQ+/5Ko4p2Ln6/1jpu0FrGjL066J3iV9tTSX7uv5tgQuZRh0Tn
XiQZKtr92Xzy9zJcWCvWlNtml4gfATntO5WYfkUhBfXsHh9g57+44KAIqkWiMI/M
hGSga2bnLwmARKvT4DiAbcjXTeCwhIEabXVGA+q1tYfIqmzHAeFySCauBfLOL4wb
NmA+t0Sn4fdZsb/FvgfITRynHnlgwbniMZUT8xML7pc1aVgjko9dIzl3l2uyC79o
oEGTnZN+LC9CUmHE0BFoAKoCHzxVM2GPoEp4oSx7v/sVZBikl8eBgfGwXotc7lds
fdJ1kKtF0J9aLtUaVGePW83i7Q7kf3jSMVE/bZgQ0x6lvaS/23bGNzoHDzyw9Y+C
KG/piGulHZf3Qe+dohb5BxV+45MTDNp9CvEUHAdHbcj18xJh1B032R7n+iP6xrAJ
nyHHIHDA5vs70GGuL2WPJz+jiD0p4LHnIzwiQen6xBSJTuUSahBC9E2E+KTCZ1Bs
T33owiCGGvfC7v2C0QvgwUxrEe26sIHOtUJDzFj4YUnLRc8GuwEsuVgaUej4w/a5
egMpNZ408vRpRsDXi7sChVzuYxQPe6iMIIFZHgv9Fu4CjJaXN1qRuaha2kv23BoI
EYpGeGzMNhoX0SF30QsIgdJB4zkYReQWqjvZng+2M7gZyAdGlC/DHJD+sJ+boWN2
0lnZhIxNFTB8vpTpAj/o9VO3kuoUPNrMN7tMuFlwL+gVpCvc2OHCdzo7xWYDviOH
BNLXwnVr/WIVz36UDY9o0/FM8o/v2WbwxmvG5w3cltTNa3FxSv4I9ZiET0C+Ca5d
RIMJrEyqprH33jCKiYA/ZkjlFiuoyIRJRmdSS4rAzbEQnaYBwd3kDARV3jdThqR1
+7XGA+cij/p8hauvajWjI+RKg+flWIuPmEVeCWpyfbR02sgUd05saHnYK7p6ZLJG
id1H6MJ5cPZfMTOe2L9/CqtfHecoxUAlAJMFRrdfh0RF6RI9EI0QMEzuD3L72ftk
Hc4U7PM/fduzGDjXloVgg2Kfw/WP9HXj50LslNAzCAQ68g4J34EfnRTZ2SFOgvaD
TbnedZA9C3Y7DjXXc+gyaSwjWnKKk4w8A3lnfZkAA936pdhJYrVM5OUlzWnpbu0w
tG/2TzHb90wMcvERkXOE49QHL6GOf3mqFnaZfLOtJYVesROcx6jRB43eh/ErKTWv
7WXyOmggeaiZD9/ZdeMKO6x4sx0ON3vL61sE0Pt/LR2tlUjrXLiQgvJ+BfEDKJDO
FJvkFysOuxSNBYmXfrhF/DAaUxrdDDWKlxnIeFWHCcSnN9N39MrR6wJTvw6jka2b
g8xCXR7zHtiTliD9sFu1yWBhhimcofzNpJmSJn1JgadICjauPsIOHBgL0eXp1sEH
ktrkGbCYrvrJFAt0I9vGOjz5LUrSADpmZp5RnS4dZRIZnltF4/Q2oJf7UOHyGscB
V6BNn7kW+qF0pXMAGUhY2gkrxhOda0N7/hRLe5RpiRUAhHZjRGk+3vvVKJ/e/a4c
ixYYhzNCRx0j9MD20IvonhQQzRK83Z3W91wQqdz4ziM9xrwbm+SbSdI1Lh9FmHWB
4GqEx5j7nWLcVuxLAujNIzcI1zqXJJxRRV3yYeuENh7CW/g/KFY8+2XKGwk2vLQR
ITC4XofDuuQNoe6W+mIyMddAhRvlB5QKZtKlEmu74hq9SOCvQSsCru/za2eo8uMx
ju20P2e6BG0HPWVMLGIXkJcjmLWo3ZZD1JbLVXaSJgqWKjis/8+C82l78gDx/hpL
2dCs12m6tNknFxvucERErprUVIhQ75o5koE35XV5EY8rQ2YHutq03hiBLFZYyjYW
wRfhM1DODYc2OM0WWWaudNVEvtKDGWu9j5zwyIz/iTBsjJocHPk3u/6th6HF03Ps
mhQyreq5xyZFFRoTeeHjXZ0MfWX8VZiIxIeYFKtzPsPhDRJtQsQVaEhcAadsheUV
TQ7C2N0o2qetyy1+WIu6XM7tqoabrSU2staA3ZNfsGdrfZCjIr9jU+OUr5M9rtcO
RnTlwrgwtedyIJo2J9Mj/2D0WSig0aEfB1OMEzhebLjUq/ylfOSMrJbIOhyazuNm
bXd5SDTqJQfKz0LMvGYwySQ4g6iNzamwmHQKOtcwDesfrIXYRxHWTabUBlI9jrhM
lQRw6SWSTdkwuIJS72ZDgYI4GtXeEdYcAi5yLYoL/ziYIKT5oXfOSYMOhnHlfDQT
P2RSO0d9INg8TIqbqHuOyAghpmT92K/ML5dLznfCfUXX9BhBePNfLeQs0R727kET
tRFjF0TnhmVSsTMFVskBfW1Tf9o/RFBAyH2dtvuT4W2ZQOEbwjAw7vaQm0gAx5dC
FuKMVjqdRv45GV4VkLAyAMAjvXRTjKihc1C6d1XQvedqEtqr0gxdfTEYailBsIr8
Kz34J7MsJCJjYcoIvaIW8eSZ0wgbCg9ivOTiQH7q1T+EAj0hEanCYx6gPhnvSgyB
1CY1L3xLdoDcikbsgIsTPuL9hdZv8F9F4CZb4eh3GcAaJS7hyZWge+JBoudfC09h
XWh0ppb3O66Zs/QKRE0HyDn57qtGosI4owdGz6MzzGZiQPmjXYboT+S7N6I6YxjM
VfMR55BYRSCatdGyFX/swUnxqNyuPAEiGqarFbnus9v1KnAuVOqVglp5uuUdDf6+
Ak/PT02x3k38qyVzwAAndfj4YIBDdY/FJbpcxr+CSEsOXjD7rnZQmBdUPUo42Ejn
EH9UAi7PfGBCxQCuaNZu9SRC4mQufcFadTPQSdR6vIcXAR2pdVqKrfUFeliw/Gpb
JCZFhOKieU6XtJlUPxizc5JKE0qIF8W+hogzGa5UjJ+xtJnPmVQPzqdgSfC0eqlX
3eEJHY9NjoaF++RcP/HG/WWzyDfZozP2Szt9wgbJ5zh4XB8U+e2jIrvDIu/axdf3
0JBpFzikxelXn8voFt0D5RAZxTUGBoLsQMLrU2gSwg53UYZaJMy4jOkXfM2Oz4bJ
L7ecp+2y288qbDB1HvUHcsqa7Ee90uouMH89iWCvkasX/lGUSQ1w6QDSUVUjMvQM
igubOpMrbsVFpGndUwB6gb6FkHin1O+S3HdggnTUpm8SXEAKYDL7bYOAD7SaOiuL
UV8LjEczRGBLEHVQrAbpj2yQwKcs3295jA2hsfVoYQfSKeIWdEuGDzPzhWGtzKh3
BdLIy8ZS9WNoW4QXt8FpUjbc1xzsmMjFAjusyHfDumJbDs0bLUVIZklokABdsV4x
mZyZg5qz9ZrhIGaPazkwMAegBH4+Cvs+O5XCYRxUOS9JylGydULCiow7PG345IkS
F0tLiOoPTUH1P19j9e4qbpCFE0qg+myVnHYYXOmr8x14Y67FNyV74QNXaWBUzxy2
8AKDsQAu8w3LUqZj/wDa3TE2OcNeOzR/+ruwtZsVKZ5sD1CoY0Xea26+S68kLdKf
Y4EwJJhSGVWaT/9i9wEnvaaIJ0Le1bd4/xzo0BmGm5aeq6m4XhAi8AxDVRfbS+4K
donNeNoq3JZkDcCooo8VmrH9OZTGV9dKR5cKuHDoortmk9JhKtvohqdq8t5LnCJx
gJ2UW5i1N/NtaTto97/lqOFf/oEi5sOeEe2hVgsMGbiFjPbnRMAgKPVDtb/Y1K24
VlZgSyX0Q3FL6Nf11iiTKfRmz7ZtoCPOOkkA9siZZ0ylGySzZtC0ZdwbRf3ezRtQ
2izleUDMkuwAhf/9T2hFPmXCishY4pDU/rYg6NPTNlptaJWJi09Rwx1omkj3HAJu
zG0LwVWfPGa9AiPOBYrNCy1XzTOJcwKf5GuyOp3o6TBAZtIcsFki0iN1c5RUYLWv
H1xxNaFTFzNDXwvS2vTjD1+v71/7cqSqaMuXlHC/1+NGd0bD0Ed6IEK5d0O8y/Ue
hulk4a7v0ECTQCYCFfCp0WRo02/0+fjoqBOzLa/cKD5zBawZ0KD3jga+t9NgIUvx
me8u2wY40LTpacQBRyxMk45udqBTXwcvL00IR6cLvVQViizIW99kcyk867Mef6/I
raDl8L9oZOB2VFn6X0cCiXJNPwxxVIyk9bAXl0yP7J3b4TW9iey+j7sTztZgLsfV
RvA9Z8Hg+OuVGQ13CI9fJO6tHLm+eESmwAqyOGaT4xeGB0oWbmoaY2xmIMXFRImJ
w6FDeGx9J65e0zIQ7x9CoJmNC3mSckKC290lHNWgHszxcXOSEmY/tERIWOkFNSn6
JosjcFkvS2fzLIW3FFKt3yfQMtBYTwmELYEbsymZa4egdq6SDKoykY4O9XkujA3k
LDb8HM7Vn2PPJ3uYsDYgaaTRfkwKic+msNL4890BRc+lG/XvDPQnNVPU1WoD7AUE
q7TMfEy+GoZ1F4krGT3IcYXLkrjm0k6bu8AU6HHd3wQuIthwu8XBV1aiS0B5B+yC
xsqD50iC8pYmZ+9BzyZturB4FyPdbBpawwRTgR0OHBqorb0fiGGIV719eBn4SDx5
k14wbzi07m/9pGetU//rWb6fE/epFeIZkkDTrEoL4HYwLawomzXBJQr3E80Sje6T
eUG9VGWUlIphORWnSYt1xGSaE9yDhIoi2mQiw9CnQVeB6YFvGz+d6x+uK5MMPJJ1
IAL3hs6Mk6NY5sHlZu4wNONzkKJFN7PSarc21CoXFC07S2pzwI/o1zyLyPEBoYeL
2gori67triHPrHm5E+VZ2E0janaSyMKCXSfCj/qE5yMZIfe/Vz0/HnSnOVGBv8r5
/USeqB2beWUPX0qDDvbucyaYeq0/NJr5npLkHoEg63BLJDcNE/NejvTIOhmvQO99
e6Ffg4Iku9WdicDj90YE8VgNfeI6a2O74pE4X+WIRrK9Y4E8R/UWK9L1/saCDYXK
2VjUzr3qiTrRLgJTMtkC9GowhcaJUEF9V304aXcI6KT3VFlbE3FLQkFZzSoD/lni
cATb+UtaQn3AnUfaV7GQ5f/p9YkPmLdUV7vYrhWPUmdWvrniKvHVC6wkXEfSJJZ2
8n5SkUNtu+eH4mjjJ/TUKoRlpAiInqCbUy2rZaRWdzjuiWkPpNkHPVO6G7OXQ2t3
ZeZ8iy/pFnwyCSM6we/huAGOquWhpXu1Y17DRNqK/p5eT/S4/RaAs1lJHxtt1xqL
fIPjdn1lC5/BvKW8Vy+1Av8a+VM35vKMjOZM6GW6rz47RM9qhY6oTHNCykfq8slp
22/KiF32oa3a9ln8uFTBdV51zyBjN6oem+GFmKGLInz8k9KEiQTNoZswKKoSk9TQ
RZSKBjpKYUKD8M8rUoein1mKqF0lQSRuI+n/7eiqpZ00swLi5O4/ZD+wEebHbGcS
nkO9DebSmTvz7caYwUsq6QO8pMFddojAMqjf7/UlceB7VsOKbBZDOQisSUNGY9jX
Tz3JjFDMcjENQAjgf5zqH7Zh/z0rIk0wLE7WsagRnJwHYsN0oFuNy91E9dQ0jVEP
/ij8Mt/cVzUxILn9loeuG7Yb9JPC4csc6BMwfqR+2oGQ/Or1IZAVTD5nH8J90ulM
erLYyVLh8D1MREfKvDrRSbpOW2seb8D08jqIRBiT2CzXlHm8ZStmhW5QyifI4rzW
MrQTJCt9tz1lWFyRhIdXr2Fgt4WNGBuoj4CNguMXbl/iNoEcZj0Vn7HKLy6CzP4R
C5i0wQmHXCuS6vmFAHMD+MPjJ4BVZEmQHwztZ/gBp/trZtNeGRG8gkKCu8cYESBC
vj6gyzWM73I1QJxZv7j+La86kvWI/mx1gPT/6d8Ja05+GGXAp4aKc7OPn958Eh0D
mkeu9MViHdT1dC+V7/SkcEshpNbaZFSzS99YZypT63rjdTQB0DKS6zrkg7AfHRqV
zLay8XT9d9e61p2hlOkIeb7VuIuPxsPWBu5PZFpeedAbyu3Co31TZd22PEo+XYNh
1+GwECJmlWQV7/pGyEr24vownonxNQHKN7XNP8tHORpJKz9+coM3/uZkGpUHE26I
5K+okilhcwMQxNJHKa85J9aQ4bvg4woKacA6rad+YEnD/PTVD1D0ErMXWMm5PHRF
EJK/jMSBnwMe6pEzZdL2khqVvX+GYOnNvk29b2vyYzI80d69E0gQ87bO7WzGQr1l
2ZynvCocakoHSqcQN8nquKfQIEMRy9FTDpmU5QZa+7pZBbm+a9vu8b7mKK/fRu5W
pl2I3OOk4Ot6YxOsQNenSbKC/RS0e//DMalbgQrufDfGvBCRxnXCIQ42OX7XGPhh
71IJcvkP16FAgVVoFUcGGUhZxs4llpk6mwkoNTJ3qtXV4jd9saCHocrRym0//b7x
NBaeX2cqLU19ZCKuG5yrBTs0R0psQjQ7E6mqcaLceLT/Bg0GUV52qA7V4/xjR8A0
8s2x9BaCuPn0m9ql0fKRrDkVRq44vCPWb4o2Kr2PZ8JJ/agpp6Q+0FH3w/1YMyCW
c4lGtIlxk2HLpaxXDmo/d8yCTBaw74DN3IVcR0uTnjoin99ZDF3014K4K1TpQLLy
/dIjVBYogz54sC2ZKg/+cuB5ZdH2YwFERGTvRUZGoCXHIo8OSiMBcdOrw++aIcFz
wMQXt2W5rOs8QvHHaNSHy/lhrkbpydAgXUvdxcZdC/AyHIImdlq+o7+Po59/0P3y
BI5xrzfjJaNxzn2wcjEX0jAIo4+sgyeOI2EypkB0pys6jPafFeqNca85uVhs4no1
vWdMXFZrVwXr/D0LdqdsNZNhdCY63oL8eWjZJb5k4+r/Wh8bSkhjTq4KmEBe/auo
Fpg38xz4oZXvECSTz7DBoGynBxi2fTTxHcz/4u05Ci8LhK0Ny2AKszpIRQSrXPEm
EtYqgEDj9WMrkO0krNLi3LMuileGSF75U0eTMAp/zfeLKXirUoCqWFboXOt/QRlM
QcQdlXntvSh+FWRC9TxvQ9omvThlImT6GTJ2Mp/0sGa1OdE2KdIEh5lXHjuzylqw
W8aMijYffWySaKESGjqJr639df5OW1DH97s/8e2x52ZjkE5dMe/JiA49CMNjXXtv
JBwfSq2MfE3EiW4bntcRDkxoKmOrWA3Hso/s4UINKy8BqDZ12fIE4WivIAmlr2eB
vAS6eevl6+W+nlfxW3pRaJnYupaI9S1MWrxFDQhCdo/HPdq0MVPLWRkeJJ8a/kIf
h0kW9PsDEHe5EV0c/qS9ducsUUVyB21dWDDbCZ7k2ALj4jiwxoWm+/DPmQweau0H
wbvPWqsaw89fzww/dfs5Vp+dSHcnedarkNihUx5aC1LxHDTB3JFcI3q4pqlErh4F
D3S4uWgf/aWDghrMssHZKy0OFiK6pqizWErFc8jx8mdOHgpsFbU6UODZhb4/7wOf
bB8r2SZ9qA8l2dksldirvqzR8ORp33i/cw7sq01nh3SjOUDUDW68q1sWDJexM/fN
6ZdHWf7T1iJHnF60eojYyJr1nZOuZFUJjNpy29ZbI6j1/aDcstyX8Ux1a8ILXuNq
mz5riaSdbRzvrkLmJ/PGXrP2RiAXzcswcEvPLQIptdYriZoPZ9GB+87r4lZ2ltRV
R1Ed+hXTTwCJoN9S6hmlAMTWjuctf4Ad17QF9D5tQ1iSZHaiLT6FvcIEt9TAvvIc
JPKiqD7SJOdqz6tIpejzZjYoECqPpiWWkwc269mgjA2/CJ+wdszOToOsI9GaHEZm
sPBQGvzDN3BLfvKqlAG0hOApOuRDb4n7tKPSJ0IEPGI0M5VMJGF6YTNQZ8/4NcWC
7JJQ76r68WtE8fH7vWhdB3OdIV2LXyyGW5LE3uqvk1uWS0Gj2LRNKIu3r3baJTfr
MQnXpgPr83m2JPbg98grazx5toYb+AdRUN/xdT9dftGNZCEBnchHwvRWuT8mNL9j
f4+6xEwOce0YhY9vaHH5MjNAfei+Te49Nbofk+kG7uYBYfmHyO7MJYSKnDj28fTr
KJ0YgqwdXO5U3lEoqDQCvXwWiUDJbHSgqwQCT7feHvy7W+IhLxAwSWkuuswtYwbM
CL4mrV5D99/7tbuTpq5cHFXum9ClANJUWvixOWq/wgTUGKXlH2zPwQXAjItm/QKV
Sdg4zsyjjRBSDEdd+UptS98l5BcUhpCqQCMm9mNlGpFbwcdQfOjr4Q3UKeMqFVit
VsnJIf7T4+XBIDSrIDeUr9eD4SbZxkD7TYSbX5oYPNvdWnmiAzgRPOBOIjbGaTrU
d0vi1skWaYH+pWQEELi7GAcEjKFkYtMgV0edQGQpSK9fq8qCBU//QhN5cUbmfcmw
TGe/NAipRPxvlqEzhZkaMbGU6BAW+64D7v0ZKPWEEyIvuvk2aE79lkxn3Cv8gsZh
l9IAggv9a4l4qlbs1Dngr2ZXJBOpaLceJcxqRMgJoXVY5iZAOmBv+eXCiA2JRvGm
2hIAPSK9MtkUf7xmtVL4s036XOnDjTIna/AqU77+81TD2H4cC5PHwvU2EFUJ4XwO
ULJpRozROLIr6yX0WdTwOW00EAsoeqtWFFlcImPZfz/DLolFzT9Ok4YLijDY5JyZ
ruVMQ1GBFHFcChZcgEqNb+ON7vSoVPMeA9gk/mWmWzVs1IMSEPoyXAZhl60wTixB
BasjexRXrPJoAEGCKWw1FkqXFulf9gMBIFai2mbBGJ+XKZ3t7zfdzTOcGHpQp2Br
9SMcjHsjsmxJERiIvgeWlnNRKRe7hDIwA9+af2FCVUbEuClRoyHreifZcCWZFigr
bKIY5UOex1fLKW7+FkdnfhlOdQ8JJov0fg/f25nEiFkrXcAEra3T21UZJ+HrhDkc
vILZMrpkFtkT+VZJrCMnH5HRPUcbgmQZG+h2NEulC8fbRywvCQHvffL8+EccNcOj
4yBW6tGuhu35U8IEBWW1GO+o2JptbXeea0yp/2Eml6RU+Xx1kcxRCMq8HobHl+bH
sjBlfiDBnNb5qK2lukxlZ+ZYSxeOHUqrv+enr/WRQTmZRA3uUAqjrd96QA1DV43j
Sl4mRK7w/B+UqQtvHGirDqtUmQEk42VSGY5WLRLA0ycrWKrKaIyLrlZiT8eFNc2y
EZ+VkEOgMJlPS/Gzg/Uj/+ObUFoVtOLTbpK87dGTtu+J2P0aVspjZvgPiw+rlqSV
I6Vz8zqJVmscxAWLZxrz1CrPTE2McUXTV+1d3KQ19uQjN/9zJrG31an7DSaVfC70
XmH3xRdoeDCBaupewddTVlJNXM0JCU/vs8VX2wy0QHIri2fOx+NaKI/WlmBBDrUc
PjjwYETVqbVJjJjHVfVxPPrpUzF/6Iqopt1JEJwrbbEeuTVJSjlQuz9SdOKhmnOs
ZvmL+Py5wDyqt3h4pPeQ+DQwgUlahaZ9+22VXuN6Wpgptbkn4HU7lGA5lFoDVlkz
Gl/CQpY70qjEnJLd76sM4oIUzt0c0wO5n/CFiDxugjJRnXjXW324gvuzH7Tcgs9a
jHwDADsjtRI7vh1fNyQcqzuPDI02TqmYchjwKgWwwvJH8CC9Uu1l6m6X+uLmMhlr
Iao2V3sHXZ6/wfmVJfnXAAwX5+qykQPzxXJcC4g36qUOPXEQMxM1cY4lVa6RqW3T
9ke4vcMcBMLsNk/zw9OUqJNmxuWgV1Fcz78eBi8uLSfwTZntLO6iGaADQQrJPXu4
h1ddzffn7grMo9yg422YHP694MxX26KSqBjmhJkgaYQG/T4N6uIOWF7O9CKRhTNG
ktSzYdr0Bqvo+cpQFTeiMfCHT7hfmwh6dFQL521UEwHGlbKRs9v2ykDwyyqjOWPX
jjSY4Y5t2zEER+cw352x1glI1IMdSoHMfUWdbpk56ezxF4BXO2H0fe0b9NYAiOEF
qYQUayFh6MoSIZ2dZnXcPq8c5xwIju2tX81BGFfM0/zr3f1sZFUC5Qv+iPkctsyg
zOu+LlPNAsZScCe29Dy18ISQqm06OnBMe1ponGQVHUkfMQLGstNzAPFIVAdTOgYm
l0/BZoQ4cCpLfbk0W8GZ6dHbHb1Jxur0uvyba9a3+bDegvBqsPcHK3LJtBF1CN/C
GFNPOuTwTFaMRsOGJuyWOZTetzboLpUbOI+z5TYqYPavrYsWeFhyAxoudNCpWQUy
qnsZk0fB5Mu+kcMnDwRdrgDbYosajublrJ+2AH/G+S8pyvg13RHCbanc24A1FUoG
xZaJwkT8fLDcz8FaErmWqaALHS9nY3givWVwQK+9OK8g5nwvDimlsP68uzBn2+YP
6vHQdRJgVIgKsF3NaRIpBA+7s2pBO9Wn8/98QtmFMHrschzxAIPcic/2dP9waC/S
ZAj4lIBKSfuVpWRrqjMOIDKaX7XIS1VBa2Z3gC8G7nJ4n9Jj+uxteUUgSaYxzV7f
LxsoFkO8aFlcOiHit3iRABJ/N6Q0RpwCZBd+cXc2VMCxMWVfNeJvv8Hmvjd7ptYq
p56psO/1RDLwPNkg1hPiLJ5us6ZUAgKQXJQZ/5rX5DyJNKcyHDbU23UUl1FJwWCM
2+OAMh3Aj1SG7DPx/xdRKyl+tM4dYpvdTfYn+/xIZzGjiRNEgsfPoEz2QUQUTHW2
pycFUrXMINQag82sExElrTDocC+NdMBjKUF9OwpWIZGKrLw+GbquOsbWIH6VKD4m
29ht18PPV9RIKs1/wxl1bs+HgtJOevBWk8hCzeGDgIKYgoEZ8VJa5WFYAZtwQiPe
DAsak/LAPFo1iFzCXXXNTRQqT2NN7U6+AgPEtqz/T0hz5btulCrpS8ZpeP6MkZfb
1coLL5imNTQ8Mt2QQIKKRvrZAEcWdkLZ5mWdxJDEMBmOmpOb9B4Ixpp1zkXWb1uB
29HTMvh+1HPiVZzDmVdoZJO3XdMsBkxLxzu0HYZ2tND6lJpVB/Iqp2FkdhCVu3w+
8h2mTZ55ILa/Pe5Ppi2EU3D43K3h5kpDyAXQw98zclqYhvdDh+NBt51TdG0OBLef
kFUwoXR+SvXsk3WFqmYR+wOq2sgCQgZgX0j38sSz7qO4S1IlT+bFJRdVhgf9LyXk
EJu/fckhevId2TQAeyb3L2IVPNi+rghKJ3Zox34WgdUQZMPnh1Oig979ozhhcKvY
SG/IoIFxgVZI6efI+YHIBnMVTLVQVDQIsd26aTAHBCXc+X2/wwlIbjHYMYvL2jho
EOk2oNh0Ukx5S2ZeYOH34qb8DXq4HJaWRIOuNGonTuK1qLU2WMXBUn6HUFNNenmG
By38nFKvh0EQlqpp74gsg+vnhHw9Bqn1xAZfbX55GqVyYnI+v+vrfSlqh4zN5FoU
WVzMo7z0EY76meFijG+yiFOJMJrMr+LXavf+yW00NXTCJPmVknMoYLvnEoO/KNr6
pIp0rC3SfwgY1ktGBQ0Q25PFr6ykIvNdSpTwjgkjH90WZ3HYN6I/7IgDFnhaH6WH
qTJhrtbjr6MHTZwnUe72hv7IYiId7pkSIlSCMLh+niC8eR9PYUiQzdXBYIYtNXua
zvqV85g3Z4qSgiblFdK/Y40bZM6Y8lW9S0C9M+thB4kVyAhjiSDreu20uuRzLzbD
DCcq/LqUBP7V3uf9HpQydThpBETMOHDZaiDTFrBNdICCsCUnIZHJgn2uqzl+O5iV
h6O9k8Mji5p9/F9DbLwZ1PEgBariTQ42j/YNPdBAXiBPUO2k6wf8S8KxA99j9Q80
l8ERbwC5dCDt+ZiNid21NcHltfQqu9orFVEJFKaOH8X2S4Q0DtRPg+wa89ayOBeH
MO9NgNMXThxTKoRQkjXcr1QKUf8BImzcGPJf7+9vrBLoHMyHrdSB3/WeSmnQL2wr
vjnox0QrxPO2NyWvK/2smp+Yd2UN/Mqg9+7Yh5Pou2aQ7uAj+1NfkcFW30Am9IkY
LFTDePkOj2K6ESbtTX+Sx8nQ/8Ne9I7PUCUBpjJR7sKuPzcihyfwCJpPOs8nDe7O
df3Y3JmJhvzImHjmbdciuFxGj2+RnoaNjGu5VEy835IuN55Hs2oOcmpo4gkJpeMm
0fA9mAYav9UywqLUNHua+btJsjpEjf/re8mAJMQO1zvhipj8gaV78dNEAR+aTVAN
k71I9GWxAtSZ8MbO+zhAMVI3qqy8XGBfMunMjiMVJfRwxHOLWFIhfFle0HR70vW7
jDhqWIbkHA5ruUvnFENCL/UL3LjZ4n1vtodqN/VLWi/uzB566NZQrNNnHkKOHi7n
hfgPnQZ+RuTJ4IR8tHP4d8kzwKEDp8qz1oiwJ92metlv0eJ69Z2vrV/bcVQ99Crl
xz54frIqv5Nuj7XGcy9ppN6nGuTGfgghASztNXUb75PAgdX2x5Zsa/xGj3A8kZHq
zz/y3mF0PNMDOW/8pnt8UFQH3sOEJBYWaX85s0OjvPRn/xBxEVq6WrqNdePLOASU
v7Mqdz/Lgqalv639vsW32R76NNfqwPJM3ksqGkMUWN4FflxJ3Lq0usXxPdr/Qk3v
v2MxKi1QBdyzUdr3DOeVRe8TzcZRReHxIdBxofFuikilwC2KaATU9O7jzOeD7ymi
jX7qNaDECSoWs6cvNvaGCJx866F12Jnu4qrRC1N4Qk2BZ2eZMo2OUQqug1O1Cm3d
vuVre195Zc3EyMiFZWmL7FgQ/enRTnUdn0wsdV2/MmEFYuh7gX0maPgTaqK7PRVF
bvtS7YF0z3saZdirtkATttijSH9fYyxNR8XpnY9KHawKdWlVa30QyXRQx1s9xbUt
QEajToTMsN5HyNpQin+v3AemgxubfX+vCvzPACdZPJnIS76ZV4AZTz2Y0B7i6Qp0
71TwqfYTFpumaUsEiiMD/SZouhAkeoOS34FgDWfOjVk83P6jXdzF4ADqVnn7x2ap
QG5OgnucUKcXPFky0HzhPXtJyzKZP3yU1ZGUfoAOfsLeTgpjVZ4xrXMTgYl9dXV2
Aso/8NgORoWZyaAXSAv+MWdzxlCMr8G7FEkH+bxNNcWxE1DnKUTmmocJ8uuObvbF
4hL5rEFpJna4AfCKrE1FjjITYuYIbjK7UMRVdNNeKe5SQVU+NbTAMrKLC2QDS+HC
ERPBrfaYi1szbGchotP2NWXld4ahnutRkvKDaE9vX3q3TRg/dKiIPlfkkoAx3xo3
WF3t4TTKOg8KmNRV+8I6hj9L8ikGZ1c3THIxP3KtMg0Ys6obFL8Ujmnoln1Om7mh
JX5YWIInO+oO4FEvCVhbFdgeHt889H4bm/twsTqZY/ugjtsE1EWWVIfpUeqrAN1S
omGdvbat/L9sAHK034E8K4ZsPjX0KupmlEOKwaUEvtKlFtULv9odQ5dH191Fml6X
KrtkjVXvL7wEJY5q3sg+R2NOmDDIBZFPRK4iAaGhKq4XS7b4hvpyCCczjn+8mZ/b
MH8xxICrCbLfDRhqbtfcrZj8oD3g9q44ZtFGp0lbERPTfleIlYo4NieIDbCzRtxb
RJBEkJk0EmdX4PoUqJzExK58DDaJZeJ+1CS7B+vhbvxTNj3OTdS3RCRQ43ervfkO
UAmKjEqiV2tezcGRKXJxnS/+tq3iEaTiSs6zfUG96H0H+B07oZZQXjP4LAyxZ8o/
ME7tWiawKz0lLUgkY2lRDu7Bfo0vxOocwqfJfv2uUdFIlBFQZeFVsW/wZVpIuuLG
+EITuUwrRjMbElZCrt2PX35NyoiLwh2tKi1dpr+v8DpZy7MhijiJMWSng+Sb0IfO
sO2wmBBH69rKcbIRGvPfAzvCqEiKOr285nIpbKLBsH0uzwmwCm4g2zU+NNx5lx+l
C4zryJ4/4lj3czVGyMmsDvg8hLQEEKcO35JKFyTMPijmthS6XqR3KV7pxQ1F6iJc
952tC173aRXT7/WS2+ciqYdfw1NGJ0jklPUR9UzIG7gg1P8q3b96Fah3PstKIGRT
MoIw/9rWlAPJivU1Jffq1NokIhUPVxO2XfahM9bhtZfNEISvXvai2fdV5hxBxuGi
awYV7ZWpqIADoVaOmz22+K7RhZ61DKcUWvBplUH5wsIVNQI8Hln/xVkEviNeNi3L
ZLlSYm5+tKF1jtOa+6t5JVgbxBJ3pcVwljKuCR3mT/RKBQdF9rcSRCEtTHOQeb0H
cjOHW0MqJOepo/08epcL0ByfbofKjLaRL/+uh5xUA/jjzUG7MSGMZwprebn1iun3
ezvdxS5I/AflIU9B3ENGwTSlGpKHL7me+1haCsiLso4z2K/k5ji+A9kSWxo5rbWf
razR2GF0BBu/yl4qeUrOl6WCR4vvNVrktEfYMd44tYkSjxW89IgBzhe7mNbnH3Mr
+sigjwMTdD9DLB01Syb9zewC6KElrWGyQi5Kz7JQaTMPK92cJJ0r4PddVVKBl1SO
RjOBL2uucQVgYTCeJe8p6IpFFEtHJpHwgXlyYBxpoZlZ4d/1pefRf5A/SskXhwe/
RCoDye9M2g1dVRET+kFOFqMK9NnebPEHmgYhJKVZE9+CB28npQFKx8RCVQOs6HQT
DI3TM1RFe5qaJHHj+n5CCg3+K0LOxcwYPgeCdNN5zeRVvUIt6KQHpaDQNZYm+vdm
FgzBuw3sJpibX3hbtkM3EZixQpHAHg2Sx+037Gh1+F1BSmkQcQF4Dg05rzt70A6D
+bzr3KTY4c7ADPH5WcS5yySzmTxRzb0/hwMFh1mw5TXipBPXFiNzEk1xlw7ALUAi
G/JA8ImCYfwgqdukO7QaAoAB0+BN/B1CAfte9c7GFuLavjzu3ow7G4l3VkOrCuu2
asJ1rVJRplLDp/JtJVNDj6ypLfqiyUFckIYh9Vhy8zNBi3xVlhoVZmVfK08gJnvf
WF326TCApJWFylvXeVbHTq3Mev2gXOPQojT9J77lJdhuNkxOntiZFfjSTcQUm/0/
t0qSXLtqzhvGj+2RKxhnmZ9lfQqBNehAoh798Rb+5pGpbCLKK2HWl7Mwsojnimw3
UWnIBztl5S+AomoZFZeHFPjMkRElWBTP0gfeo2ViqQt5ZAnStnMuSG5UIb5X+a6A
KKZJdtWUR0hkJLU8yCTEB8K+4YqITyO5mNMQm1pCyF5qHU7nx8lI9XmPdd7gUaZ6
2UXlaOoxCq2Xw5Qc9vnNOnxgxGb7QJVS7jJUFHulClYKyyQ5LO2sDIJmGEEIipNX
n80257lb7k6Uv24ANCDJ5B0ldK6/OIxk64p0SkbRlGTmMdF9l7SxvfwjfF9J8Ond
omFfyPCO4UkJ6IsWhyMd9YZfmG4FBFQ4vrd4OWEX7gR/aYAmsQ8ncNk22rMfudvQ
7vF4hv5OdjUAP473jYzJOtPoVOTV7fh/3U7H7ILZLZUgUZuKUza6EQbEYWyH35me
wfhCv/gsoW9pWeI74wxiDF97cWcicpbedIGFtl8+njVk0liAjImVNvVgl5BKQnvZ
tSPzFfVb+TcjZMqZP7oJP3xA3odxDzNOUjdFCj5RujMz31oH9/woBLCRsMKyAA+b
YIAPz4TDyRScJClZGDV8OtLKQ830nr7Go867+WzNUyKRpupYAlEerNxrcEvRKJXs
g1CYsZ/JTLUImIEsd5Ux6vLjAwlK+8huomsCW//NnS82BB0jMo9FYAmpZxqgxhGJ
mmz95gTw97Ek+1SUsOBQyWuteUx0xY0aPx5V2VBzqIi5JPHq7u1PzCRQrl3FKM0M
sCukR0DAcIsDCmLSVDTHfc9gaSzFDnSVJtanbaQjZZaRQiU6J+ToLg23wdb2lSXE
EI6jCHftBacx+/6IxjmYuCJ5kvoPbEZnmcnpHYgYKlwhnE16jXweRaJEB+IFYcLH
PuPh5WpnosqzB5/xWLcV+9QS4NF83xcimfg5n8nX/5L01SZaIzLBto92Wy6RRuQf
3ElWngCLflC5u2F6Kql7Gt9sZ783H/BeGqDVCCx+4VyZ1806m7npdQKE9pnc4xxc
kQU1bu4xmAi7qkMSMS1mNlQaLwvFBW1Op/iM/M+2BKZwzpvvOO+aQEm5XRSNiyiR
0OVMfme1TPjzFRwEbThISZk1NztxxuwjsZ2BA84tZaXSk8kQS27rAURe+y+KkRLa
GHPXzKnSpstU8aLwPvlK0Lmu5goQp5vSIguguGA3zGGr/BZ1BXz3CkoOFnWwF6Oi
4OQEWHsFph5QvzBxkgvHeqMJ2tdoEV40hffbfoPlO+2Tj7HDP+fPzsGu6eHMXca/
qFjBbBG+iZn8+P5OE6yTpm4FfV9Bfb7fEiW7jyHY0UAjYhG04as3kDEExHHGGrpt
H1IxNiLhunfJpm8stx9akACkJyMjYMXFz1IVhSIoHAtro24cgMHHJW/obsrQW/Hu
cj38DSrvEpV1ARDhXtnkOYFCQRFo5Qm6eyjXHv2TepPDwPzlf1vUjaDOtfPeqqNF
134hVIVc1TR/i4Gb1Kiz7gJyxljUGDWg2XlqntJ23OGB8guj9HEhnSLhfhMKs8iJ
SUIgj4uflinlNg1LA4++iV2jjtkUxpWZueouo4LLO4WGNAYv/KoARp7b8Y+IZ2hx
5szsgEFYq2B5tUxAwnsP2Wel4reWoJ31AUMBg3TeBp1mj7Sun5PvdgR+br1765j7
8UsNuU+AoRuZ/vQ6hAq/nrilpdCcQihgD0Lm0oD76A7gUQ/KMrBY/9H/wivBwjdo
8A+myy9DWHpzf0n83rayuicVlQipWQi7R1PH7GT+fZ/7GTUREeUbrflWStB2INNJ
iVVTlGluNTCbE3SSRRqkcvH2rYE8PLS3mVlWqfZa6seRoyzhT5hjnGRXEVIHNC6b
oAG3aF6gR7kygJEZii92Nqt7Y3DSlfXrMXt0BtYz3Ranx6+DQJ3HEsRfehCDJ/dI
TNzvUOoOPlD3DP1eCsuEEsu2KQgC93rx6RYiz8mnyQe69Eq376NxiE3DRG1dSvKq
Tm7namsLkXPRvFJzSwaK353JODDQ06fQB5HCuc5A9z4xAl50JdXZZnA3aQVhAgMu
tNQ85VCrzIyTT1V07/1QVFoRX/BCCmuD3u4ttG+qcgxswzjEPuTIuxvz409keRxH
Tv64/u665dlTbvLAudxw+pNb3MWg8uvFKxGtlX8bMGXDraAwWRxJaCwD8JG3blaN
T9Rm85Ky9BOfhzhEF9jm9z3YqOzWKBJMXmQrEyQwa9p98phcy8OsO4HLwnPyEneG
X/2hPs+kKaE8dGUw2K3uqGQYDpe6JT/6J9aVkR30W5aW8Fue6s7rVg2FbQcXRDW1
dj2ebKo3iXW1cUTZ2rWL89a2XFxBbAv3Rw8jVzrHNnCKzh1Emzzpb4u3177C4LFb
2QPS8dVkwcKZIyAnyzg+gbCCPmmb+ehTmLaLzwp03mZarHUKaEWOdojP7D/oy3jM
aFOir/QVDw6dB229eNPyyvWjMFrCjk2wQzhHvvPZyJqLdI/VAQaQrFkS+qvDYdqU
Ts6++9F3uVpJ7UTvllIMHfnaXsBqHRISbmfKxE1y2ajbVZAAsEMooPZPoEbj8fuq
FO+qQCMyKxlaNkCIftwQDy4RxVTfGk04mAwHnqWl1Yn207+vcTiaJVTiMci4/1hH
BMfPVfMNveVI16LsRd7BjXjM+gEfkf+MD0U2dOnzdcksTPL1cCclGVPrSCFXCzTy
c/p3XbekVxBdbw6KJ7YQu+8VZAQpMlmCsnRs00FTlh7ASp+wabCrnFCa7kq0D0Ai
sV8MjJWGcJgo3vXV50nQsSv5EahLjQ+AM7fw2vbBUFkNWG4gfQwEVQb+wKcxzFDF
QhB0VmGRbHCwHB4h4Vr9BQMUkDUeTWnf5hZKrKdRYU+AjLFcnSjVtbw2YOtAu4/J
zxxaoP2+JAHO+I4M3HP6iZ0SCaZiLSMLhdV/wdUXh+GIbS7VD/Iup+rk8W7PPNKz
VuX54J8Pmr0N0ikFpjBn7ZkOZ2J/NaixkzSGFmXrKT+62xMefRrJaPj8P5EyeRci
WIsxC2yZZwekgPCtUBexxkLSyPKOwVSfNgejlc35AsP9rbVdY/646diHp+AKGXfD
buddq8APo33k+bW7ljkcKnCnbmOSgVxLeanE6R3TTxcrWlffhYhNXr+/+n6bQcqo
DP3Ta638sKqaWkyAJUO6A0QBw2BrW1Sobm+U5Yac/VwtaC12x2eiz/W3uU+rDaXD
cd1lDwlAJ0ru4zE07ujG7DyCJYU3Rruq6yQshrZ+Cr/tSIxjQn2E6Oqa9vGPyHkw
FFB5iWwY3+ema0MSvFY4Wq2uwCbdg4Dle4okzQtsnorGJ7KsaxzDIybwiyRhrcjt
jJbVtaEy5SBkOK1I7ZTyucFh6NxoWie7zjaUZgELbx0c0oCBpWdaE7tjh3ffqUgr
UdfmI7cc/xNCRR/7dbVK/RQ8CLKtK0hqKqo+zo185AJXPmcbdM7flzPgFk/PpN/z
3j8RK8POkGamOktPfdS3DTW+bCqj5tnxsaNsTFmJ0VO2HHECXXVgtiPW01Y9ppTP
J2+MpVP7Deitnb5XMtevY4xNOH0UY5LAAFxvEtW8mIxMFiZLcYGwroBwzE5e/XfL
Ds32Zd8NkzEZDGMT5xzwAGTeubzBQwBFyGra6ALMs5IMUzgZosWhC+6rm4R1DOFZ
saRG+ndWRVqLf1gJv6btfW5z7hssd4VYxx7ExMmlMCahwTj55tM1uyS19UgZ25W1
i45r16fRAv4AEUQLwKhjGenK8h6Eg+rN2W7ahUBMEi55FmZUUhnPDzg/Y9qpemKs
h7Z6R18iUsMTyStf4oo5M7k3ZZoAdyIjAVlC+zH/z2QE8ovAP6vSnVg4v8OEkGHR
FqYhOdMOeXs6NIIBk/5k8p8LpI16gzJuU+auLW9sNSla/4uhzcOzayntMn2zIiaG
n3VO8PELNXpLmlgAGRrChvMkgvXiDWrMgf3MrVJ0s/leSCWUU9Ayf54IxHrKuxxK
z0kuAQ03k4CtWndb0CFBe+7EqjdE/qXCMD7S8HwB16N0a5HVFs/QSQOXOHM2WB7v
msj+DjjiyaQw61Rv1xOQc7XWbamzAWHkr72u9iu5QwG6b+rvaopvo16YnAPLf4cK
MZ9XAFMLX8oypC0k/99TdaZ4zKLkEd8R6h8LUCOsDhp+UW03GP/v0QulPqroz0CP
0E7smP/TAB1YGoePweMoGmbRFhQnv1EFHBsRIyrjA+iPai7vfNEU9U9gBhy0Zf9R
5fqcaD2or7DgyYxOvs5xGqYDEcRiKfrNAOad4CnOy4NYEVlYia2r0ZyomMpW8CPf
NhCrVBIF5lyM6qysXtKhoFZGJpkVJhn3p2ta+b6VNxHWmOJoVO/SXM1cT6fahIiE
v4lHoOt1pKe7OTwfscYut0OO3bYx6+iwlrfKflwVIAiJIYSbaFk+u5GF/JzCLXH7
mTzCHmpzQ8NgDHR+aKtp6zZ2MwFZqzDke8iq4jbRWEaUSyruxUJz3N9JxBnewXbj
u+3Zm9yjBNHdDrX+kcUoqKyOzGTO5jTV9Zl+PCa+ANfnuKdT4bSXpoYCKtP+hH2z
7oJRx1WDlvK5W3ERs2l2BaA+Gza/WFEzTPFexqNOVwVk/YAzKz9uv5d4381kJcL3
advnVqmVsTYsQhuvi1Lqijo6ihu4QrDUvuWOWJSC3vZDqV6Yi5CQTlZDHTahpK2u
zM6KoqL4pOZvLiaz4oxrhvDb3HT74oy4qn289kJ2LwEWKgrLD9IHIv677AHRG6KE
2APcomXEPB0UfH4yGtSCJNsWz8d3x8YWuB75xd+AFWxCu5hUR+a+2sohqKlVLQgC
TTlG5ePPCTBwzEVlBK19qiKCF1LwW8P2ugTja/JeJugBQn3xJOJHgrsrS+fesUsP
bx5602TWys2uR9eT3lSiapMBdS/d2jQkXNDXen/BSzY9kGP6EIKlS09Ce7TszmiL
EKeXj2QB44Vk5RK/8t/8gLF4MTHIzYl47fE+2DbJmp4MvpTx47Ja32ezjaz+KQ6I
UpS2m4q4iBYxHzrKMUR4ZkUOX6v01ppQMgX4yRuCT3lqNLwqf0hiZS43Hz6hLMLr
XDz9YFr5zIZp2DbdfmA/jZF6bKh9QoyC2860tllx8oIed/VaTuayU10M0oJhhcmw
hfdpHV1igTVVO267gtXCD9Paxo2pb1y7Pko91lvEsGnSpiEoIyei2sDtHH9M+IYx
piJnk4fvmzZxhndJ29tjrxMlqlBVp8rlMp6ZNwQjVgYlINf0rL4DeQT8mbiyr1Ix
TMjY3j+BcL4DYneNwVcBOY5TPT7Wa7ZgBL02S2UPR+oZJBX8Hfd+aSBi6fE9doNA
T8QIPdcNaOAFyYraDRfNmjm7Xb2SK8os3dlNjpVpylSggKTDRVbMJh9LEt28XWLk
4maFgniTXxwb8M5d2PeEyRhub1s5BX8mbFJj9kdlha7t1Drn6LjD+JplR506EeSK
PfEiDOne0xt63OnlgJHE7TCapq4FO3YNel0iOb9eeS31cMKbnqJ0S2vCj4sBSVqN
GdS0jwhCnQXnZPyll5gqD5hDq4OT55Ka0xKIWOYsUrb0oQD/Zow5D25jTiTntGXR
NGz0rX1FxGYrMIipBPfNim1g1RPwlTgodSTFNjILmzkfhwjs5PoIopIXRTNc1nwc
H0PVHjPc6vbbI3jvUg5JM5vY2FkSTKH5q3eJnVXLJ2cLWBq/Z8Cszlj0IEjFHmh2
tgzTNcsq8sx9SHcUbb9POKu8klnx2hoMood6togjDBO2KvLML0Kf+ebDHYkhXDF8
BFwy/KOr28bBglnFSgZUnnVLn8TeJObPkZl6EVoJP3n0YyTcwciOTdLbBS3X1JpY
OeAnAvWBL/xze+N148kzeGFOdUqYqbUx8ufVAmH+t1vYY1JsVt9wRBRsSpZ65pLq
Oyt2wXJC5ohP9mG15PLhyLqoruRsR4rKnXXPLH5TKmSifo1dADAVj1H0vHp4N1zY
B8NEy7bXC+rGcRp3lNXcZvCPq76tdESu8m/0OI06EeWmiBGqcAyIoExfHwFZfID1
2gcKzQ77f1qb+/YW8T+Fpsx14OV7Dbt7738WBJSxjo+kba8kqSSwnUOkEjgs+4Ps
YlRGdPCy+xU9BHc2HZPw/iEoD2jdRDmwOlSwSKlWuMQvCd8c39+++17skiHwwaLs
56wnlz8v0bdzl/Aw4RXevrTXqejI+FF1cikWljQHv2Qzy+SjV8daRN8BmZPI9nQZ
Uk8x3PakR/nn5o44GaTXfc2AWdPv9ZpDf3Nev/XC8T0ntXZ9SNEHh4T57t9DGUzj
/NSFDGL5SGJryqfhwD//uwAKYFoIl+9a578mT1UvAiR963DrIfraW9RsbFUkhp8b
lm0CRdVM103fCmVZdsljL95EvTMTfQddwOGIEljZMbvkjOwEJ/Za+L9NEI8EFNT1
Jjd8ML+NXb+oa9JXixqiCBR2GMi0MbwIvF7Fg3bZHGeI7pEqBZoyhmO9AxbbDg0O
q9RjwjuCd1v3Yfq0SiG6QQZJRqbU04OUZGXhVIGvbDu5b7u7kJ2OqfxKdswmtVwh
82wdc4m63aQ+sN9nl3OoAnYRAKIJhRbBN591tVxdcOMkpSfiGaLLbsCTg9PKoxCF
BUQzlppvboYWKcCbLdvTN+Ubm6LREWofcC0CTDzCyCNQupeXMw3Z/hVujFKejZiI
O6MeNF6QCYgul9l43AVMac6SsxFsZAz3LEgzoI0pfFQNZbLc+kBPXic7vUL75QiW
GNlT0bh6aDCYzsBJ6z2WGDWCrUHT7V84sz+8u34V8L6Z5eZicbphJH/PtEOBqmjv
n0cKT7yuY50b2IL9I0j8VlA852f6t493Ha8XEZQ7b3cBfA6OpaYCCJawKyBGohD7
F/Bp9yx4eDCZAerl8LkLZUd5Qngte2Q+E6878AmZIsCfgEvPiMsAc4DOek9o/ZjG
WMo5WAMZ1x6J8Swpb1jGWOZF2DY/fQ5Da1CqTEYOY3eGwSOXEtaTnxErPdKTFBhT
xJ/LdVmXvs73jcosIf6C9ezBmJHnpcT8jOSLzkWz1I4qwGpDPFH+Ai/WYmfcspZx
t0gkWIRl1WwnpQaFKhaPmoo9cPE40HbPDtXLU+DeDzKolytCz/sTsWK/9F4txVld
aqkK73KYqZQHNlsONz2GAGar8+zZUtmmiVxBZH59eawOLhQZ0KeCKKQNv4Nec281
F6Qsr4U6VKAMtKglTCbh2IbD33wm8cag4Q7wbAiVY3X6nKY8s3Abfz+W8Fj9lG+9
jy3Nkm5reOf3GU1MQ3sIdRMb1LQLwWdcmGDqOXzdnqCYIVWADiEiG5HCq8P61asm
d1PgiWPmwbzdXw1v7vxq/QF8otlCfFOUqJ+EbyxXqZS2fFDbwyJQf5E3jGBxynOr
6UtcMSTWYyn+52LKAsx+mi6VZnie+j5Lw0uJHAILZ0rbAhf/5y1tSY4B6It/qL7Z
IcD4w6ZCdwc1hEOAS9gmElluzOqDZpuDeoeJbx6q9J+oNQ1vF1ziikE9mLSLG2Ub
rDAV7sW6n653Seu4GT2FYAGfaOVaWnz1+aXMfJ0Ov+YXZ6d393hFjjtM2obor+KA
OahVtX03xNVQgBX95JGoTRPayLK4QjZ24nbkTtWuaKZs0sO8zZ+z5dSjx0R/pICE
tOf1c6iu1DyBRdO8EqwmNuxeV50qvpYL9D8t8WI+ST+OGoKkLJhJtWwf1j/q0EJD
yS27gpYVa88X66LzjjxOJYRYOg70bmRVFm2xZawXadLjUEem+dX5GGZp2iPOj5Fi
N3uDS20yhp2RaDwj9L3tmKRuW4/bS3onSuYGrnRaffC6VV9JrNnhX035Z5KPj8fH
1PQucYBuH1NTxbfBeMCyQFVxewPf7OZgcyDPsZfy2LiyOc0CrnCkMWKww7GYBivM
AiK3o6ucUc69cflKxpR2KZUvsw31ZBEQ+xy7q7BNw2IQGsfExDZTEkS4Vng1wip6
LUbRq553/RleQIP6CDxYJR0uSgHoHoKIrKHWXktgIFFsZYavCheDy3kptRbGnXQI
a9g4+I8PyccE/o8veeNTcZ8UXtdXJAkCrtZvYYGbWJM7SF0S1zhmtaGslPWPJ/Hf
bNMXrrB4fFDhOtWkEkWS+FkwPhLBUQN0ibF1lO7gnYYHHs5WZV+8K1dGneLZi6e2
dnABB2eq5dZT852trQkofcymo5Kxeb6Hy6ANpvxOt/rtQ9zR20Dx1+1lJH9SlDqA
957xsOce897BrN3L7VYMxNoqABUOCsbhuYM7huXa9QN9iNyc/23NG0q2oLnOSoqN
QMWEsEK2uGjObjyTobDMNWdLp3ffnCLVO4qfU6pnGUlntY4K7bJnfd3ojHVygJte
Gz9nkuM+RM6igbqhHBHwgg7hp6ACqqZ/UVPxOMDATZaBnOaDaoOJj2iK8WSFhIPD
2cHwWPHeVCmdx4JC9a3mlZlqib0dktt11o5NITAySX0VGb900x8g4u9htoJQ5xPV
eY7MP20q/3OgFpS+1m4W9e69ZEUNvHIVGhaF2bNX0RwpEcHWCITHW9BZHFnpbBLV
Z9nsWnMI9l/32gkvxbSXA/wc6WwEYRja5B3KKD7aHRZJyLyDksAQqPJ5ClblanCm
yVQsdgxIOMmXxLZ5+13oqw7GJL+FWNzQjJ48zwX5DRGSLYIShq9aZDbeMTOxKQqt
OTJwG90d6DU8h1K4kYf42C/jf0iCuw40R+2hXZCHSydLThhdj5vwsAz+yymgi0Qz
gYKxI0U5Qf0gye+csUGR3NJ1yFvHhYuEeLqPKC44MkCC4JkOhukDcGKOTevyBaQb
MkBQQKeZlYAQ40aULn+ik1h1lCYX7uslUPT5dVNhQaF8q/ySeO+rkswkLN631RXn
cxTXl92qwHqX0FiRSXulAmEHBxMt+cUsSMPPAGUTKIpxzIQ5HwtbsIrnb8DacIwf
uRIY0tKA8JL5REGSpU1dWZD37135e1isi9kS19dVpN0o43CPrw0S11lDX31NbyCu
re2ObOplAcKXFrQ128IoFEOkqek0LAudhaWWrEMT723/zZlCNybqcQbkRF/p7z/M
1NUDcvNVbz6CvS+IHoKZ9uZYAlsqgnHan9zqebUDbi4yjFqhsyPR4Ofe61I35L+k
FWiNovLdHrXTULQbCSi4fCuvZArJejFbclhnnNhMuLIvzKfS7BiJuDNBLaFRlEPt
PtcUifFR9fTwQuuzxczFsuPM5JRNHZ+GtJL/bRh5iNNzWNk736TbFqS9Q1nI9NeP
od9seZvaVYErjkwQf+OsZmThiwjIp91jGraT81Y0jK0/ueZhkstmdqRMGYEH2ox2
HnrWX7+cWJ8b0XL6XH3CGG+eXP5D/Vepp67MbbSDmujr2K1KFiAxA/Z3CX0pjaQ2
r3PhZDJ0MK8f1wFzelwSci2w0YtWLQAUmTgzV/Yu9FV3k8ELOvZ3aJ5EmkP38Be4
qZ33Qohf2V2yrngBa6fgnHg1pV4BZHAD5/rblx+lem4BUSSihEaVl/ZYABJONjV4
Y0qBeY8JDrClAsUVcTdKv5sTiOw+PnAzKmnh5JhvZrftWBq22iARnSXjPvh49xZV
xBh+neMKrm1bmh1bh9UrkrXF8ledASIAMDT1K/2kg7gO4e1JEfui7wQ1uZDTKq1G
FcM/WUw+PWf8VMb6Tu/pjN0CASzsYa9t6lpnOhKWCYLUWw9yc6u3D5BRRecfdjqL
uYaB2VG15eEOq84KMYDG0qBHVOH2baN2cdgWM3939x7e1+1KHqGLJ2wys1OrfY2u
MF1Qlomw0Bodw1Gi02SaB2b9t3wcVYOdgStgzTGe2OS3+hAhNcq+Gsd2xxY/hkLq
K1Y/JI/uElHEEFKYUsHBBxXuudFbHqpSOpSuAX2TS8+0uyRlzlmQu/b7S9b/H1pq
U34kfl3P9Pr9gcxQts4DNqeAdajo2Havs4N4aVh2EDeYhUoIcsVnoT24q7MTMWlR
mSGctHxY/9Ws4duMvgIpixjHGuMliMbOP5dnZs3bjY19/o71rPZRYWbbNMD2r4ml
Bxh9fIXys18vjW8FG/JA6V/3CqsVWZ8Jia9UHk89yGMfiFSFMB+nTN5/HGrAZP33
pOjdGsG4GigM12MF8heutrdvTw/YLgQpoJNOZrM1NWDj+hZkKs2FF+qnAwhPq0jQ
aVCY+cQbggdqNi0A9fGpk/l8ebX9Dl/4CqgNzC3IoBz8mueE/Hjbvq6tYBgl7ksn
wvU90S9fsUOrYxueBc0lnR9y0s7ym8sQXOc+2MAvUBFuYtIZdz06yYdYM7JuUmhx
Gt5YK0R5STvJzCHzbjdDGmH/+WyTTcmUFkILlgLw5GJ/BlItpgadmTFUm6DkT/eU
1OR1sKqhWPw+SM/aUxxK9tXwm5CgWej26qE0K1gABQplSiVIk8HHlVXt/w64Hvo1
BvMdAl9bzOUiL2Ks++/Rkoi+OI3d70YKKz9ltwF4NysuN+JAstNGDGmn7fo3V6DB
oTZ8dw4VKzXaZOQW0Z4dvJe2FUA7+XrhVUKnD9v3QQzLspfBQKJgWeIeiTjbW6nK
YxpT82Gh7L7iAZ3MJqnu0NS6Yo2i8ehofte0NbfY2+XRF8xJkEirUTlO4zFFbjjm
4yYYUrzpKHcxP2syTmA6TNtN0BoJu/x53+qIxdbAcVL5iYo8z0tohvZudIepk7I/
eVWvyNwLx3DjavFrfNvFxgAZ7fQRLdmS+1FwYYm+y90lpnGuvovAjw3kVdQ3bxNs
/3kiT/PE4NJxSwYf64U3uDXw79JW+QXXIQt4tixoOrkGCG2GFtQs4hIG86jYM5wp
GZ7LRCMvC+XdKvGot0XLdNcKTcfWkY6owKmkf5/XjWtSn7lZ73uXPcAO3jGsfhFi
Vi2jRUn+tHbtuRFIy3gGAyjS4ZpHufnwbHOU2sIQ8jqxdlZ6LKRk02W20qepRtRm
zb85B+h2q9k1cYiVhFOblUJ/MkiDFXSSWi9vWkQaq+FDI5bXzo1ZvcYaF8wRhNuA
nh6J3yq7facQEnGmYmKK7vSia0GsRTqgXuub8Cyx7ZKrAjUFnU7ye5DGmQ07RGnr
2PMCmO+Ng7tLZqsgEwlI1BaAfKa3Z7z1bPzQwlUfXIlOk4mgLqljivJJJoof3cEm
/t5jTLlBptVZqUd8EHxQjQO4I3XXs/Iol0agmNhkEGIcgbSrPyd3B2CZQpsUyLQZ
ktIENi8PqgHRnZ2/b4Ry0SYZ/rPTRwjWB2X/82Um2qH+1z+UggJLtGx0ZJ7Gq0gn
2tRFx3RiCSS82SpmDgMaeh9C66VU66fC4YHadrVeGCW6N/IZ8Hw5AuyMEF4wEjsE
sz+t75o7RxEfzoQfQCb2WuweQqyRKO3jZ/sSJum5p32XovTzNmrStsc1OQzSh+qu
k2K5cmTHdT1vr4L8Xsse9Oyeb1bWAvZLDPHTQ00dzxR+hyAhg0FgNbvxZllzRSqe
HKflPZyRZfbtwT6CMtltpRa6quco/u2tr2N2v4XGRDdngwrRq7Ld9H+PbqjmDdGc
Pc+f2wVAxA3KLvmY8UHSzdvTh2Oov7P1ZiFzr6IbstM1G7FcngVSiJAXNqyGXpZy
/DmeGggqbgJorTG/R3FwfDs6LbFs1U75lYVN6jfhQ+hIWTrVH7e5pWQqccjGlDUN
OQ61EO/csCDZu6dVY9d3HoxOToYb9U9SvZ0KTg8x6hqaRyH6Gd5fy/qNT9YliOJR
xFTRyMRnvKOO4pJ/X+zNyYZ2PlO3PszFWukqRfRKu6yCg/nS/por7yQYa7rAJE2l
ZCdoZyAhCGxiP7WB115iQXLHHrblEJ2dCBgupfZVNCNilKIHSBeRGHMaLJo2Aqdf
wkwqBC3JvtuDRzTc7QEn/J2iw6Ug1qjo7TZIyQoV2+1oWzIU2HrH5Cqx0Gqzt5Df
931Ej4Uc+S/SEvneYayw2zwYiIWzKX+658kTVI7pyZRC70ibSXPa8HdDZM+8fvst
/aBAiC2YgVgrl48eBST7hCFsSHlDGG7aY61lqZgrWuEyAUuNtaJ/4Uob0CBNKiyB
Cj3U9VuQqsKSbteNFAGcO6t1E0fE5u8gZcJY17hq8CLACVw4ITJ18t/kO5AmZEXT
WQUAmjzTiKm6+B655JmhS83SON6wQlpBhO9P1cUhQw4uW3EtO36tV3SKDf0E8p+f
7GzBjrXEQH5xPPdamvY6PY4rrM7OFkqjSlH4IlCa+5fVAU/ndA4MentxZQcODuOi
Z/lOdoKWIgHo9vc7zbef5BF4JansJ97Fr9SbKzYuaaKO/m/NPEEvv0dmV9tPYn8/
YnWGTWqdsuB1fLuVT0Jz39+MtpOUX9SPjRfRuUJ/zqfyGLFeX82WrkR2uB0il5ZM
aqShQJ9X3FXnU/GJtYErdwggk0Kw/08UteFJDkShqTUUKZhPNE0IOwfy1WFJcK8p
nT3pF8rll2MsdTgkm5OwNuRAfmju2dIsKma8SNUL6bvnJOzx54ygMXLcdFpnNg19
t1Wqfq+pVoMeKRkV3wfuPnD2wLxjDpPfX/RaQ6JzpDTzQZthV1QxC7rqLOTxO3nS
jLGHaYPryWg5XZHHj8C7Ti4a7jyJ0BWD7P0TUw+6uvGwr3aXP2K+SRwTDuVxDqdG
kay5WEhNvQGlgtnc7A3jgBts4gMRLEmd5vRJewvh+9AW65TSLRn9qE29/2ch2Mtg
oB9Wvk+zVUUJGV/VMcLTtVY1VriVl+voapdyDZH0yT/L68m6wUJ+HiTR6AaabJU2
EKFVfJL5MyOR6d+SXfiWVCiUVr77OzNyJ8SWSwsEsrP6FvxUJf4GPdY0ymo9cv7R
RDekLUQmXhMQUMlYboLIN089aBIaH8Lx4Ew96PthEtPL/7KpDM0jozJdhM72dsX3
tHtWJfyCAJqO/H6QeqXxk9tms7WNydB4Hrax8GnTMs8KjtEJL/9iryiMV04PddrN
BK9QdvaZz9LPvb0hwWVz3Pe/qUk2NqsnM3HJUsyUWJjwC95pQDltuvBXyzxWGXdX
i41AagvM6uacb10h+uSMZVI2525xgOgnJVI2kP9Xqy+jcXPILq+wJe8awuY0IOVx
VZN2I6GFJMw+VRNMXLladGUJvsN34X/5sErRPDZNfswOLDzGAatloUih4XSXLQtL
5/avavckpW94MLb5+UkeQja1atW8VzcvyUh7BGEjNqH1In7EK51IuPVUT5IHqd/T
sNZe+9zppucBYc92KOICcbpcd5jLCceiD04ohK4ciM/WP2UNHCf+b/mQbxa3QH+f
acW0l+Gytz2ccuhT2vXEl2p4es4qcX11ymGWzJVFjZgBaykztz+CeqLAJUxdwpge
N42mpW/Y4Co5We81o5Aw7SuVH1oCTMjfwkgcqumk+Mm+4sjHHw/y1HwnR/iCZBWA
Tc4A6FiD9AJuBbpbGAGewkvXZCeI0Vp60UcJ2FZOZx3bLeRvuAQUSBcKUG1EjHZ1
m3uhj9/0940ezTpAFasKyVi30bnavZnlv3q4ZUfiT7wmIrC35hsvNM+yPPzCPZiz
vBc36EWRnyvKKtrelIQfO3IjDliJztJRHeuBShSJf2LwCoxpSD3dEFsjdcs1uwuy
S2jmi5m0VpLgJtTFpsQ2cffDSgUpTHvio7d+uPplIshVLgJNnU3OPCuGhcU96P+Z
CF9vzD5vXSZLYsJSF7U+Pj0rdkyqNP+HTNH03B9e97U6cj4LEzp4Nr9urkrCOkcI
c5NbFLw5JNk5AUIKx5HqW0MVg8wcXCuTprVdo/Auhca4ziu29touPQss87CqcneM
xw9EVM09hoRMEld38sm7iqRCpTWqdYSMM9F1Fwi6s9PO4ERDY5s6I4urho/x1fCn
h2ZMXMQuJX33D09iHP/QS5aZveWte9w33JSzNoA8UrLar/qUbMTcHOrJfa+agMFe
Fa6hpaKx9xHGQ7U1hMgCfVJzB1ebLdUOiyM3KgDSqdjT7Em6/k7Ea4vZKtjgCerg
zaYe55enhdkGf+JiON862EQgE5oUX5i6hzyV7tcpvrD6FrRExRcJ6iVP5+8TApaQ
QZ3H0ug7NsJK7S4LzqZ1RV0BzGqk5vxDrngegPeHJnemz7jztzZqQT+N9Ez5E9uF
d3mpfAe59nczsx3d0wGzUbD3/9PETXYaTTrC1EHUvJCwupa8hCZdP/Gk14oOjVte
xShJgD2QSsShsZ1xmBTEsMVHltZGb4w6WT2w6F12997VvvnV+ZoziUn3lV1Hg2iY
OIKyF6zUQlAmenmBjDm81GRH3BXXplUIbIIfJVoltblMXVAeE6yt1p/ZlE2tgzyg
+5pvcQeGvvPV1ioK5BKCcBdjCsdqvmNB9LVBAaFK5NEo8SMp2TcpY3uJNQhFyjX4
7Ijaj+ULG6BrRnjZyA+cDJQy/u8nsK6WXvLIeYyx3WsAJe8SOXMVQfqoi5Nd7QKn
Y4P53HqqqQybX09ZdlNdcysJImcHXoo4Xzawd1eP51EIMCeI3RoZmqnNWPfhRpwQ
uHcTkoMK+A5V/1LH17QdgiAfrpU4epyigyYoOzkHcJp2Dxmjd7uuMmzrLgT+LoG6
FhSW+9srNeq8+sczNF3zousx3ChFh3JAcBn9920zjJg/91c49UYYPDEnfMn3GSl8
X/UchiEEg7/ZXnfMU7omlklPI7yXP1qUCWoGHlhplchkKs4SPP7wTFmKSi1kPC+0
qR8p8aPJ9HgO6XjEoFrCOm0A6U6dLIe/TvXYEmooxiU7saYhJgtalYbnKwP/NYTI
QyIz4/ppxXjX1i2Y1bCL6t4DO4ItAFpz6GSvBU1rMY7s+UbrAk5Xy/bQCIFS2tgx
3isBp1B/QK2gu1wM3mFamCnVarLXSqW++i1Nx6ujWmjIIXBJjhHY/49ZDFTzW9m2
ABH2XMC+3y7BvT6HjdM0aQIhfKKuBGmMSee0cV8S+bZGSEG6/TqjjZkh+5IaTU/p
zeIn0oO+rSrBGp/1oGtjtH3VaghySW1lP+f245SbG6TNFz3vTurbTigwwuuVj6yX
JJce6JUwcwpsLSow/NlrRjnBrfS9W5tnUTo31wb0/jfzuIPxvELCoZUU4ZGDvlXn
9gfGdt5qrkFpjIdLjGaQHbUOkNYIiNK068mgEBpD3/HCbcHLATwPw/IIwf/3PKLD
6enLDLILGNw+TQI7YfReWr1jgcrB0YyBWJQvYpG/3MDtsS6VJNgIqffK/sIro3JI
6Ap2+TkD9vjiokbblMQ2E73NhXPllLjjrSO8abXUsp2sfsu8o/ebZRDPdkMHWNi4
ScKWRuBQaWgts/crKSQyeqJzUt82zk/zZpHxx8rUZjt2EJv+0unJx2rcmCjx6JS9
z43Cb1DTS0MftObkO7hDjGRfmAgkLKFyKWPTKyVD2RVPs+MU1e1D8kVujlmG0hLZ
U4MeuAOeyJsB1DuriG1XhMo6ln4AEnUrTbklL15/WQVIjoFkSy8n4EElSNvLZdIT
8e4c09QL66d9gH8MNyfwFjWt3uPHUiiTuCbNXRw2utf1uaPWmgJaImdyhO6QmA4K
x/deoQMVAuInYp3uL4qgQUmXIy0wQSfYuGebrW+c0JkRcrkblSNLeKqalJkmwLmy
ifO3cQp98FE3B1z7bEvbUHpvxiYGUQRhZoDeidao7YtyFLmaZJkvYfK5Q87Pu8qC
t9qWqz33nXRfBxakL0ODGPsKhFq5oNBt/BIAZYyL+D/TSCbOjG0vtLmqn7wDZKZt
jjerEbPh4sW56CSGEuYbWDl5pWFhyjBRCUEe725pi3tPCsp6KgAGx5wX+n8+Fonw
hMMaN1Jn1dP/7CT85qP39NBZw9t2CPSIezyFYuH8XzbPSaR2Dj/RGCsN3E1JiB0t
GY7tcMCt7JkrSFKvUV70J1ynJnUuYV+IhIVP9KD6k07P6kWbB+Y92aM4tBUOnR49
Yw84iywcuo4ej1j/1jftY4MLgnkYu4ZTqvmbFa5z2azdJ/g5ER73W6FZSlurDJ6Y
ShEjnjoKtYvpnfHFW5mQ7XuDC3lZvggYOQDW+04/Q5atTP2+JJ1iZUj0/bGY0dLS
QgYbztuPnqQVvQJtXeetD/WJx9HpkwzQzwJzFpc3UG6Mfm693JsJuqWGMBzn5vN8
VXWspJnp4hn6a4mM96VN4fit9iDETP1ECgtVqMOECulWayxIONRa0DAgCd641EC0
NzEKzB7L7qczlFFTB6CULCd/WOa2BCSm+7HIPsNHuI8q/fCwngmjtKLvWV9BGXiS
dR4odSL9dD83h2RbXiUpE8OzzW0XNobIh2C8PTAE3QquDdLLGEIiA4YajaPRQU6z
gRQbpeRakm76XmZNCppyvEDeKvg3MLzEodAYbW1S7m/0NKK1EhB6rC77nN+H8Ift
z4myuRGIBhJ+QUDPoGNGk6LwTFfZ4kfZBRwAeXbwq6g1oCqU/L5hEC5UBACU5KmB
b1RCui/KJIv/VGRbFfI4cQELQh8QKv8WF6n7EkVZGKvVJy6NKWlm1wyDo6AYDceB
v4VrqdqeskKtQQssd5NtIuxTEW9ww/JfIltLhPHLXZZ4Y2/06NYNctgh77H/EF4R
r9Yhq4zz0uw0W3v/DizhgzcFc47k2CMbOZ9bybiAYfWmlCCxgoZLcgMyuoBabill
XOLEOL4I7SnOYSHtwvAeMR7cRZkoGO5Z3rLDBByjZezfpxdKt/ock/rIFoIudb9N
Ym5KaS0rSXUl+0rNkkMjugCYjaqAjeVFi1O4DCIxvv655M3X2yr1bx+q8uKaSX+I
1Yua3RlJgBFlsnYtWBTHBNy+BXOHFydG38m6za2Sjo6iBZzYR8wwCrI22FwQMpd0
z6E4VH8nxNEMgrbi1PFtffXoa0Ijj9O1rDT7xrsW2WNVhK8EQ963cg5XyTO1qXmM
S9vlU4ex1T+CSGBK/MoNW4PVCxcIcv1hQV0PDaSlTyk+Sktzo/WbNOHOMYceEG5p
VAGhAYFKjvuRgkbtY7HwKFnZypnPTeBdKLbablRsBjZJBzbGbIsaBvlVtemnIO9a
2E5u4KT6qO/mKLqq8uLYpkWw3lz89YlcOkOGRxSdhxU4TDblAK525vNkBVvEOu/C
i8q4CiQZipfXk5fUNnPSr5wzrZBUk0E/WnJWPkBhGEYAyOK6giEtbPE8Yeufcqhn
pk7Odfw/0PsoFRU317sZsoZc2GlPUAWef7lnghygGiQjnClExCTwHUqKp21n4coB
PdtjJiQRgeIGuCxk7ZD9sOiextODFnIapPi4KhFDv7+HjwmswK3HBb2fKvBIndYB
HuMqEE6+oAgfLb6b0hmbkrseLMsoAEaLGpAVtrZxP0NePRugQMr3hifY5dLWYR4T
N5ywr56++U9wkf7Qram75wtuzaz7Tya2maUegvquBW+Se0bERg/KYHxRup6ikGuk
NUkW9nDgermjBAEEA8TD9EaOBKbEMjntWsD7aPqTsimCIqu44lE73TG4KBNag9Y5
iIfAhzYDDzjd8nBZe+m4wyOdciS0iCACjFo6/nMS38XM6yqMdJZE0FgVDy2zUfod
I8+jRTo6eTY5enJ4IXYeQNhPIbaUXRyb5mQTi9pDhi15d2y1dkMue01FLR3e+WFk
Ox3g1zD53aycJC4whvYoGhTQG1cDVnahBiZYk4Jv6PRX+iE8qaoxy2NBpGEyp1Jt
QV4sM9WnZZMf+myipx6Yb4dFK4FCmgPEybK4l59zC5vffAvcb/rvQRjO13+6Piec
7hMyvbhKdbAgbmJDdMg/2GIyuQtQPGQEJ/t/xHVaOlF+DAjB6ZoQOTI3w9zcO5+f
kfVXwBCZjBYUl3zXR/7dM4YLECiqIBV7vDpW+A0lIV2xkkM56HwWH0izdw/R8zO8
RTbkukyS6rAvuOTkpbjjoNDGuEd/dE/D9GKPjR1o4nRSOR1E22XELo/9Zy6wkLoj
3tBU3Pbe+85ZETbQ/RBqn8oZ5O851zJKJ7pBEPvawqB0Yo76ruOHEPoLZUiB4KHx
glBIGppXh1OkBwnxlATvVg1SB4mRodYzVJff6FBd8KIp3H3mecnuiNXMJK1b+emt
nqHKLETNz9yoKNZQE3Bo81ixFoIKYNhJRTvr/WhTqtCorFXS3WIqOB1leryPIBsw
8xmgjCiB6G2eFqNdn5wvbvMVnctZo8uBaHmOdiZ5k7oWS6SQH5AyWjTzby40qD7c
Iyxo0UUMiHOVU2NEn3nAUM/GZSsiyP1ZGhsbFA/8tqr+PRj2eIVoiEnVDzo9KCoG
fYV7lBN/6ZYMA5x7IjTY4ju7mSQdH11q/e/xzLpMhLsMcjCE3ObHjRwpbrewmAuz
wGP8hD/p3KsOsFBsqgjsm5qu7iIIhrAt0EE0tZihkOVClSmwgZrt4HXsvfBP1PSD
FP4oLiq5E7xNypmwCiJtkqa9EFYfe/WTPWRvXmclcJv2HjwZKORhm4j4TL2fiWa4
1kT8LvAFDnuYkUK9ZLLNM64MdbqZuKyIt6q0f2D7uqoMvTjgpzGZlDFxJ++FvxEh
obi1XvC6I4xCGtYRuYGTzYS/bZTNXwM1kkb0bgCuFtTbl3uaIaEK8LrIGS3OpHxb
fiDkaNPIIFQrFcdUtJOZwmFI36q2Q1nKEpw/r16pFQVycOrrMYHxhnRdUIuRi9/0
L1NSfZ8w7mMNFgLinmeODEaqdtfr2i2Z5Ift7+oeacqy2CjHay9MSeWo+KaLjjoe
nH+hYcco7mrzltf/owsz7sJPNV+p36VCrdqbbFS6j18C0PjZzQUDZhOhB8MXo5nb
UlK/2AWyOd1EzXV2PLlrrxU4wY38k/06DUarVKhWsaamzDnr9ALg+1Tlf2cX4UYt
tc0sOICeU6cb//Ef7BSST/5OgAcCR12BC+R6IJuo8g6ktD49qXoFZ16pYkLa3GgJ
2QODOBX3uFTgOGle/hYByg78lXeJ/rKW44mm5KMBykKMVU2Agx0nVC63E22rHtDN
iN4oT76vj8dKYyDwiHof36+UWk2CFq2EtPnbvRD2SLscDk11v6XFK7v7bXy0F3jf
V/8TnTSVHNv+ANfMM6mc4Vzsksi0rmcnRYgBFZL1FcnjmvzfTiU/T15yyfOios/y
qC1/u3iJYbzSUD7269USBPV0YeAi2FCFChK410vBJmiySU566pHv7unzt1mV/8bW
6tUd2qlmtyyK97cLj/fA4W69R54HXe+C6+eV81HWiVC+3n08JXE1T7d+pMzoJsSA
XZS3sVvVRtBZJRCTkR+8mhS8UOLIYbqdub0/ugKHYpEPNCZzxiO7i4kcamh7gL7i
Pm3q1WKy5MvYjcNNHWr7kFXI0I85ope1yj7v+0Dg0s6SO40D5TYKUJLB4c1L5lvM
bybv56yG1VRLMnnXIMvZYtyg/Hy9iOxeSBv3Jw2eG4bbdDuGvcdZ0GkwPRyLOqZK
buMVXttSqrQVPBFsVvBNgTy0Xiq8/wG6bNrOUsPqXNS971m5KeWd1/gwjsQeM+pr
xBwrtKfka9vPbMqa3qvZrbwXZqVABJHiL0iVKFKLcjojIlKEZ/KVKQHVvVxZqXEs
NNdEoyoVWOXog7fld+6VqeBRxOhz/flNgS+WeAkQ+UpUfU8GCBE9btrFL/1aXWif
d/31RwzeTThGg+PApCmFTt85/B+rXvYHk6nULhw+kf8+Lvf/Mzue/7i5Jrln6zjA
R4EFQE6aqO3ohG2qDZvUiNMDxvr7H+l9jbNZxzx3pFkDvyZAgiuypXnud0fIZe0A
k/JIuIVCxLcYbdcLO/3isIsIqS7xZ/ASTwH8i2ojyvEuc0DCnAdV9/VW0WUxJh0l
M5qIky0eQclxarlMzj7UZOiiCd5QUJ9ZDr9uEPYkfDnJZRlAJobF+begJXYlkNv+
ld4rC1GxejLtZg776ubSP2KdDGXTzo1YO08ZefUa9EPVPXqm+M7mDF8f3rmFoI4Y
MX7ZizCU91F3SKGu+myYt1vwAfW12iS++OUSwZydNYmd3pYFzjTbwwI/1MZExQsS
I09tAm39EA6UWB7/iIvMBZ92Vb85jWIjRvjPW7/4Lo34a1FfafSMFX3krug77ctH
QD8z05JHAnL9VUOP4CqX7gPYVJTT9TjyfJez6aaDvRAwihp+BXuWv491bNac5td+
JvG13wOOuxiDBoDtUvfLiShvwN/XsuHD6qaQy2yXeL3IdYZd+Gp2SqIKBFX9LWWt
t7Bq8X9hZAlh/RmSWPvd2ixvP6/VtF5U83QfOe3lp/NDWrCzitYBvc6uPy9s0SYw
fb8hKrrN84Jd+QIeH5LBiFZ5tpDsAs2NEC2UWERA3PLOi3i/IaNKHlKzs0PbIc5U
hiTgY6pgMC0lpF+YqOFRUeNnyRZef/MKw2hbBS6iLAYPWtgXN5CC3QxQd82FMEkc
Id3ByBQAAaWqrQJP5rkGu05ZxLUQw5CCkOKmMkSTIiJvynR7dSroLBKIWOhH7rWB
gU5yP5XLXcntYvW98b/MHvge/OtjyzgFO0p9zdGMe/84+VKGWc0ZaCLSpccBuQdt
E9k8FOXoDqJJE0J23q4aQXB3WfIR/RrWAcg7EShaJfMWUtD5oq120+gmTfwxcIjH
z0WcI8s6vLRpKeZCe0xA9Axp3Tp3LFWItUWCpftGFPEON6Do3cdlz5e9uk0l4uhz
`protect end_protected
