`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
oMncyyWd9VuMptAzz5MjHlwUFGNUg5aVzN+v87815T+ilmNhgVdBJPCoflO1s/cc
+NK6cLHNtwdt0tpknp6PMg3fBIdwJI8kUUefmx9UnjCQ3INgFdHhd85XShaRd8o0
BNRyalPLPoZ79sAMvMR2j3Lx+WL1LfczDxi9OVDx+MveJ5jOPDodtZt1QvmCl5ku
rQmvzXn49U8bdsws3g30+7K1HMU0BQAKJxI82wECpCkzVByKi7M7U+DsUUpc1z6u
PpWb4mr/vHkUuow3vIHeBiIMi+o0MCW6wVA7VDYaQWB8aQPt8UGlwf7wHdgBBhGK
7sXH4e5d3e011X4ifhyxKg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kGZ7+pFc+grK4LO4cCHn2j4WCojbX+eRmEOI9X1k/j0m1E7mcIBA8OjJiOOlI+d9
JJPxZUQ2F2b0I0DLoFSBPVqcyTmV9dX9jmLe8923MKdpozULOHg9A19Eg8VmdehC
z7TEnvY7PFBEg9nmRCyBj1YeUSyBssGg4nCetwMPqH8=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 112544 )
`protect data_block
4aFiAQNE1VIT4biLfcBWbBvkAmTiD+0QKtbZK4uo2j7+nHPKOAYb6TrU5/69JDZG
pcRbhQmJFLZHeMr2MDwkPRv5re/SkCsRf774JCxZl6rANM8WUJ64u/jrIszOskIG
XN8FEuS840hDL4PsMsfUNpal1ggMKs+66BYctRn8ytHp4ac8DP2NNWoSaSUP/9sg
rRPioJbA81PPbZpLnmHDrFcM7McpACL8U8wAeWHdGmKwcrEH1eWZyHEGkMgeRQcz
+ofZXZA0LzUGQVS7ImGUhIfs9Si5/ZrLRBGfXLBVKwDYfcQZglBew1yQOVmPyXQb
HkccTGMESh1Y1g8vWru1FfjtmRlCXTRDcR63KyyegDD+J+KHwgcOC74m2RAue0KL
Aa3ILgB6p6MjmiEV433I2vf+nsfQEGYihH37A5T74Nqv2z0EZ+WBbYbxCIWp96EL
vdd8p1vhwq6670Jz+fV98QtLo/iVxs9A0mNgs1DVhpxplnxtW+gQHTiTnvs9EFqW
mg3z4WtFTdWaKHIM3j+/Hy2b4vOABJpEirLyk2O2YlXOSMAsWZD/BeMqPA5gcK6R
+CBh9Qo0lFc41U8xWxoArMfhR3waSnCWoTBLD/DLKfp33b2b6HQiuNClW28xjTdi
TthZ36Jen+zIH9wPD/iZ2gdUaoYhLjYOMhR47eM/Aq1sNPEPS/hdUdYaB0MUMW7B
p8WMd4+HKgZM8HmDIVTFzX3tHmBFzttbi64xcNVCkXz9z8th3Z6JskmjYST40QTH
7Yvxc2FwqoBg1GXk67oxa8Jhz/gADbhI/Zyplkwvt+FI+P1EEXqvZYtFqcpY3Dc/
1JJQxrERlEluBOFB2qb858BKWE4vVLS5qGJd4QoW3UYMknoLP52ZBpRrATDuTTDa
xNo4ErSN14ExZ9ZOCllR7G1gUF/JKbKCP+WU+87af/b64EU3C0mUuHytBvYc2KM1
KF2MwfzT9qGQn0oy2Vo+pmgUwAjg0JHaTnTFGdPmcoPUbCM+X9x7kY3x1/bmfQi6
sHG1Mwky3AXhe6u3rYeteXkydBHS7bmzghOx5jlpruzGZehj2PaYGNnZydoqoAf6
BEAVg16bd0ab5VqfVF1LaGukUECADpmwtbGijPWQzsBR1tFwkLx9IQs0UKiBM9eS
ChtuwJPT39Y1VqGxPn6/NYZaNdGn8JfCYrEJiSDP5boJ5Ff9acT4oZny0vWxnXZa
09RIzJrSRhobKj/Vovx1F0HKmQ+YAuokmn2oLl7zgeaEAxOTSnFHJyGri+iPrHMk
1D+wHsovCEV+V5CY1yoflC4nAhyk/BzQr0NwOLgs87zkcgLwodmtXry4bOxlzHdj
I9uEWEPJhW4j1tGLjbC9uK2JyjcIWPaiQVJu1SrT4EbBDqFhjWcaXFWQiBrLniPx
5GAN+VRfudZsXGkHfPOcVVuDvxFA2kyRXqDFjNMswbMND8lTZYhte90Bu42PurzW
G57eEDGy5VtMlzzX0Y5ba9dC/uj41AHUGFAwSmT/GPifYUbS4iV+40IABIxGAp+E
LAm+ioR3pKNgots+gdPepbk4Gwd0QrrT+PeY5sIyCHlGxKVxcYrr4WHgbTqXNPcz
7IMN1QzUYsHOCg+c5Jjlzj3fKrwc+VJ3AmLZ7+nXbb7qfrLYMUMENxptQYnQoH2k
0ZORwDKMiu8ifAUw7dwVMGyoy9lzA8ucdhtk+oYyIfwS2WU5qGLYcdEwhOaaoh3W
Ni8g5dhhtcChl5IgbwJ2V1gfW4Beg6u20XmNRa2XHhtSJRKDyFTRFGYYlCcTKem5
pxWbKKhwX+b7M3LktnKmbLWE5nWKdoMMziU4osS1cA6sk5DPlZZW4JGnqs6ezzna
MNqzJ5nUbfBBKZFuzx7m8+Q6zlAc5HXrDoRMwB/iQlUWvzob8jXzUUQWOUAlr+MZ
Ss+UbjIEeAo3WVIwgOyC5o3wHEGaz5/PWGqWPdjSeYna3kig4VImTWHT+pOZaowx
qtV9TUURb4t8s4ZACUGIL6dcp2kibf/YiBSoAT+0zX/LJwv/nX4yOkxf/hERu+lG
LKwgM1LVcnHIc+GG5+Y/FmqNE/WhZ1xZB3JiguY/uiij6XU/6nJWZ9/RwZTT1oFv
LUWSzmWr2KGbsExUxfhPBCnDukbWxfEDnssVPidTX6F3bwR2kBA51KboH1vGAVfW
VcVjdGPESPFHMaNJ8qzjGOgXu24wFdFDdf2Z0iLepsNToTHuG5I35SYHEMOYnzaZ
CDnlaMgHb7+yW1U/6XgKqx1OUw01vNE8rBxVkqQ26VM3FYZBMdq2ghld5svL7R57
g5gW68ScS/YVAHCjI+tMfSA2NAvCyLUhmvs2fuyO0hcPw/uMtQOgV3mh0gqsIrnq
nf/UtyM4oobgFoIoa9VSkwBqQ9NfknMd2aDwxS/4ssf7XGZUEFfS248h3xvAHk4u
QfyrDxR7NvouC9S9hRFBAjtiJL8+FjPat+ybVlH4rC9PkPbuaaHXPOGdVwa7DKqu
x6UC7ivjuhdjtFWw5sDME34xq6f+OSXVSPlfXg3rLFdag6WXSwsucB87SYhgEClV
fmmS0r7qTJwP1RgPD+Obtmv4nSLYV3iHCskkugtnBgQY1YPHYZ/+eH5/sXGP3pcW
bUW7xZsVHp30BnAs9/J5ttl/oJoSGKCwYHpRsvYECRrXDr7zsMtZ+rqb8YZ1tJdL
QTXdU1P20ghEHGzTrDsqv6yLdoKEva/SbYi5tzkwCpO6EiNLU3MsGZVWpqEwgAeG
tE9RvXYaYfoQYWfKlMge5B2qO3rmqhQu/xl81gb1d6B6e2U+izaZsfHANUdCEGhK
nrA87uRL3Aiq3rzrqo4V0bZ0QXExkOVwm/xbH8jeSORnvJXUcIxlqyvmt/Qgtvp+
QFIoxmeNVDLftZlS6189C2TSbvLFavP4PsRf7+juRfPnj624odT2QHCir0L+WEo0
Zi6MqhBgFLdKON+E26M5uPPtACoqNVqpQSbR5UJCtUmA13FI5uwFqph3XgCP2mEV
fyouagDbi1rp5HBsGYUFliUzGEk+BSKS2yW1REnNoYT/rYu9c+rIgnHTkqscgDQE
CNIztCIkL8PHrpNxRXJswcZI2ZIN3vWZ+ZShKcnL64YBv2RBUNubjHZbt4pMfflj
BdB39SI1zqsi8ER5v7koeggg/KznHCm3nR4NPgq5S96bHeP7/SUfCd/PycjXz9Sk
s8qtA7FzeLLeC9g5J8A71tlAR0yVk9OQg0HOg8ypda6qLxLTdZnct+yKSjKhziXx
p8TJhfaPFiZq7vrzIq4w6iO6jP39iz3H68/0342GgtkWsB5gHBAlNPM6ylY+FJ5D
nWl22I0CFXFIuFa1/C4Aoz17uVnvS1iKHc2sk/t6/CvAj/aViCFggEXSPO5FpZZl
0HGdIqqzDD9VoSJsHnKzqN1bdwPItWXkiLMilQcKvY2ktDogDbaHmIf6ZChHSxSi
auVBYJ9/A1DCQWKDBEpHXEYqcOTv6DvtBKjjWVkqoB7rzXPS9+erHysk/QSt2Vyh
HkN+BJoRf5jhtws5oGDTAOQYXu1unlHsanpaZ29BsO2IhB/8ctdR0qN7ivXJcVBH
fUSFvJF4E6L7EgrPD0dAJpmGJmSC6Dbxx1Fq2y63RVDUdzQOhDPjE7aWm/Eo6vBA
gB/gOM8238a1b29OPHA6LjRaTAqTQ4NLDKydOtSG/kYGYwM7K+b5i+Sf3iAZRCYT
sCJJGaf5Bhqp2pJvrt8/6julGw8j2GQLlb9wr0XDULHtFRvO0diwYurZMXAQRZMg
Kt7/IIRQhqpseImoQGDF5hVg4mYUpu7J5Pecv3IlUipa/XxWO30nMJn/OjsS/dvY
NpslcipPyEiU/eQjsoH6G2X+UQlMD6s0RIkBfEbxI9lmSR9StnfQDI7aRzIQah1A
DaowSQ1aa7T+YO7afaA16dO+5snsebZKA7eLWaaK5z6IHlREzrm2s213GBTysc8U
2Wigis3CptW06mQuk9IFDX0uV0o07gEL0lpx5t9X2OR8tVdWJWhGGMbZUywNomgT
4yHRS+o+WS96btYpG+gT6wwbCPI+ow3AieIeEUXLFHb/iCxp9DdoelsjaZjI6MIi
TSpgvVDGuGxxUH566KCu4tn6YaLgmwYVmcSslAIJdTvGAnnkq5gu6jGC3NbqAZhw
Blq+kzyVIjrlQ8Z6xSoS7cpgAwF28lJfn4BeWKRbWdoIfiKi9b0xVY1y/rnOZdmW
9QLmEziyGVL4R0p+YRjkOetDBCZ+tSuL5+1/8vpidJhdaPsFgPR0dXtmQ9P3j0BU
VJLCjnX1FlR06+CjhaqODb8osD9+52dAAIR8ZwkW+wWKdFldlAUIu71h6Nyyq8/m
s63tQWrVyWJa21vPFLXa/3VRzh1u9J1fVJPPj2rjmHusEG+xM+m2O6wVLisWVmBa
cvI/qMUmTV9MpndYX2Z1nObq2OZMttroJuzAxVC4xkqshkP/DNqZiQ5zLjTNUbjF
NJATAPTgO/WaKxQDLqAQM6aP2T6/B3+fWK0/lzvAzCAg62vYGqLyS4KbtLdk5dD9
tWMyEiT/thK4U64IJE67lwen5PjZeljZPidt9KpnLmFzLV4Kv97Fzmf30PudlRT7
0916EPKoRDiMz6HHDPGmMqfbqOueCtQpszluUIS2jd8e0hf34sHK/Xo16D0t2zBN
yNEqGvR4B/h95m9st8UN5gxTG/9TMMW6o/RG/cQG65a6rHscAEgXoowmyrJSaLQH
oSF2g+Xs78R5R6UFwzEMWCt14ILNYUevzANmbbJszoKGE9ejuetlBWUg8yxUaLn/
SXxRKW0M6iYBuGfHwvCtvpP5SDbL8uM8jKfw5g3jlroJPma5bdBUk+lfI9TZFzJG
LUvRnK/IuOn/oWxRTlKCRvkYn0S+RKmdhFpIycSdY2Oi/5zBCJIpzD23DSNk+wYg
hNrubkumMDACl+ND76sbf3sblDTd0SmELCz5n1LY3QS93TqCgkr6JaQ/Xph5OHch
W5BucPtx+PHqore2hF/eB2oQEbCWLBkV8Rjs9VJPDOvSHLShkMDYIl+EMUHiArDK
/6pdIPAIzr9eyI/5zGCYpQLc2Q1pKBWJtFzRLe73b8N5p7BniREfKGNQC6kuLDl3
nlReJc+HNlV16X6pXTs8Vk3D7SNBrqupFS5PgC7eEAMHK+m+HH9qHHaUqCZa0ixV
IHA5/uyj4Jb2wGn9T++gO7SRtfxs+ac7QUUDmK8JkZviezVmxgrjQEwmVvXuyiJW
FaJ7oYMAJowHxdfQg1tedGB+Fj5qwlU7mDHAfYFrm/p74V9lMiyI3yZw5u0y3HiJ
EzXsxkWBkOoQlZ9m2lYhkCBmQzGr7DKvKWJsX/BvdxWSG8tBcwfig73aeyBQ3g9y
Aq8Jn64EJVTEAX/vEbervlB0c9LzXO/tPuMwRGg1SINFd6L894dc6StM5Cz8BHww
Q/GQ9XAFraUN6rOExVon0kGE9VPz/Z2LCL//Oj59fjsA3P9uH3LTxQOMM3iCyDt3
l7dsLDQ4YoanxtgMSGiso3uhkSzigSHrZqUrR+E54GKrMjFBQx4oBi/MQc+c1Bzt
zcON9kX7HLCcTvd5h0uK6BY/Gk3PrfAcHZ23lBT2kM7H2qZBAGMdOn9Tx/6zp3Iq
3LBU2kq9Re4k0TrNckHeu/E51ykEXn7rx6ZC7s+RJxzDNy7d1eCYcfOCD5jky++O
7KPBG7YYIOL6L9UbsHhY9/WPPdjjUcu96eluopfXEAQY+dHg6NKIzVKZ6G8lohOG
RfSiDfKzMtoDjwd9WoxQDNd7Fme8Gh99tIk0Y1JK0dhQyXC394HeeljpYpScDPDi
IA3HAhB/bc1gUwQE8lyg1qR0CzCQeCRUdWKalPVLEu/Hh2mrMUF3Shwp2F8zJdYN
pqOS5qnqYMi7f/gCKArwAGF9YkZnbR7G96HiS3Tc+CGoOcSQqlC49ApKwt0Ux5gy
IN+ZmQ2DQVge7N+PWS/wA2Nf7W1KpyZWM9YHnTJxtNMOg7aJ1BMtSDBjsXpr77Cs
F65T5GcBcilHOr8WazgJgaTdn29LOoQ8m4TmYpzdJJUivQH27QhwxSXE4rjuHkim
JeyQ5Ep9Tiqv0503laPMhRxdgzofL8Rr/1Sv2aP/vXXf1ReNkTJWnr8E62+2VEv8
NVqgGHfD+aheplWyGkgg91NEEp6is9XESowXBNKuiDaE/8989WGaDs9xVpOJb0u9
EPPCj9fDvm1uxyD5NqJB4uiREIVfwSsIJpnDiyYaWWHNeV92aVF7EoSkYDJGqjGv
n7qtXwT/m2WEiQKL9XC169Z7pn8aItTlJ8qqkWIEzjxWT8bhnBt8H30MPPv5HpyW
A4X59zJByEkHP+vfWfWjkZXTAHTEE5d0LtNpTzT1YDknF8PI/7RcMeauIm9WL9fz
qVTCrQmOmfYZlglIR/HTwOG3+1FJZa+C2itjLUwMBnLLroyf6CG8bgoH2DfqAot/
iaJIDd7Nez1dLvXsTQSGFkIrqQ0pseJgPM5Vgg9S/3wZHP17dyjOj5HMuMmIjAWT
xzblayIcmnYEq013/yOW0KLRmDBMAy+GeHJxkruzhWWdpAzZ6x+C1ddorcaWM9Hm
siNit8V12a7oemyhXP+GX36iisSVjRcvW74cu4x9IU/hDXV/yQM3sLMll4eGF36m
15+mk3UElaS9Ple+zTP41aFdFF9Cz0gIuUAMdnDaauoWWavpS3XIuDsuh6ZqEsCx
+WdCCUe7uZF9AsxxA7Lkp93NQgWifT5Prx7hV+xhRJfeVvm3pvEy/Z8yh/kP+H9t
4B1SX5l/2jSCCttqu9L9hZCPIj53x6tFJxJ67nGWM1aWDOaa8iRRzIApaLghNabE
uCYWIVghZ04JceZJV74otE39Yhschn9UuzsEdyuPo6BnqWdPHWCAT2ENr88NlC8X
6gknwjqN/Bs3Q+Lcl8B9/jgH7dNKE5Y6tKwExYXRE34ozVgfETe2VTmNDnEe9fLC
3fD5qkWarruGq2QaIp8+cRCjKV7jCZJS4xZrMhdtlshkp8avQn6xmNOdhD/pIM6F
0mGj1FokSOvQ19WXB3rA45NkZBjy1ouI54JtnoGoLzAf7FVzqnt9VticSelW8SP2
AKQgJcSsTaEt/3B7cvWkwKItMalepjzow5JvSjepYhceBk73ybLdV7Wyw3Zex53z
rAyM2pFOeVTU3HOiBYRHupPZGNkM8E0WA4lGR2io+YUrtKgrRKi+s9++ZW7/lMxK
T7ma00DyNrlLXJTucE/dXnuo1XAWHUSUusLi4creEUMhoYXeRitz3tV59VFZmYX1
Gnon15UTX6sdNtcCTcpU/HkaEvvvZ0+w4IvAv2dX6ljRLGBhSgvCgj3RBpdqTHj1
aQVRwgH0PFJZZ9w060HGeG4OBPiTFEmDfFDiN0evvKoYEXCIdG9jNLjvZgKkxi6t
/HePdeizX/eDJL4OhSrDKv+YHO08T6is3L/TEplyX1GAd4qsBL7EOXWZnJtQ4Bbw
kpRmeh6cBf5z3TO1vQgaGm2YDChtK+RzRIRcSNgKebuoCc9PziQsQEhWyBPBVQjo
LkYQg8VSmEcWlHT1fuc6n0DFjngp1Mziufag5kc3Z9ZBzraDKD90kDSWEh8toFjc
OxNuzEG7qY49sRWn+oh96a1YoX5AS58fNEuwt/BIfynwxDamo/0DnKbVa4BgaKyY
cXiYQv050ocwzIIxQuQGLy2dxLuHcHHoTU7UYquyZJ5SFxzg4HLcUfx9LE8zzMyW
2zYNk3leA4o1vfyWEkzBPQ8DeLAS+a7d+5ULKoX79xplgpt+3i5C6hsNABL2P14Q
bvxuo1hSBvos1tsaDu9gR1ING2R9S/EYB3w4vAZ2EJ5Jh8gfZ+CuTsXvUlaDRYi/
CDySb6bbw2K8V9lMuGglUWtyWrkL7agMlMfrjx/WvJQJxRDUc1S+a5KHpfduIUme
vXJi90TNgJ3dNTvkkivG9urmX/7thbJvqcIqku6XLAiyWHLNWAptsPlvHTqdhkLj
hhb+AzuuoIBjZYQRk4/ot3QhlfPTTbNHJdy7IHv6+mOKLxc/WdY8bO+3U2TugMHI
NOsQGJBS8+M+wVTkCh014fKs5dVYfhLostSP/hvUGmwsVErXkIRJz4nWEbdQc2ey
opkBbYJ/KqoQPOrNo0g0+eJdnIrvOkt0izYGHOKD8RIl/7mDgcdaQSF0ygoq1328
jpcpmKDAAfJmZwfYEfaaKDqpxcuEJVw6FKkgf33vi0YdC36HARpPtqp8sMGKisfS
lHt61Qm4bjQMusH8fjkM42+94X7OLCVw/wKezp3QgJLa+NvyXEVUUnXBPo0z0jlG
soN4/wpS8uOtCvdwxHDo+AoX/bO+yIcrV6bGgEGzrN8+72QgqIntBhpBFg7zZVs1
KkoDNyMciLkubrq3hWBalUonGMrulKn9DgfriTUptVFTGFGTaZP3LP6ylaIRrQQp
LHlVbukYMM+1jMtR8sxeeq9VvvADkT4Huzg5Rv+LBy1QtVFk1m0KQ6k12jyiSCYd
duoO3upWVqDU8YZoPPgZUt7cs3gtmbJCTNlhq9YyR3f1sisx71eTkA4x1a0M0RhT
5OwKfxRCmKIEGfgmwWMNwSOTLwesZGpQ52pGBtGQ101mMxYum6pMhIgGURS6x9Jr
qzKdzCc3XrlSESm/s2vYevaaXG8BdIcw22koh1TM2YodnJnl7OsfTdMNhjE5/UNf
/G66BiGKrj7ihOXRCXD8+uKdWOdPrG7L5+x7+NvDtboxEvmQqTFwG8gGnsuWAlSa
YU/IL1QoJweHzSrZcW+pIH485b5LviIxQWIHPRv/zyjO0Sjykj/zl9tPo70uevYQ
akp9L2/TuGKCmTCl8cvJ2jeXzOLfyYzfRYGdqblfAotuBbf1JL5u9nPzAIoLHxj8
ZyKK5lJkmeEc1Ffmvn3K3YBCMQhMHCaQ87NM5SEdnA1uKlbkP4WhuBzN7NjCkEQS
f7KtoHI4NOw3+rcrbSYWXSnpH6x4VRNw7/x+5pFge3D/xB+GyKxlonp9EB0QriM2
JJQQk806Q1n0y+3hK2C4oJ51lE8bG+lscIzy4kk8ByW5CtpcjtfMZeSTsSwJdReT
3pchDTCwG/axLOWL2DRHWqrZQAd4ZSu+R15vaKTstbPdO1VqhRXIeVv8Xc+T4b0p
ieynWsqhbS0Dv0jOBHhavzXZXFzOwuwO7CX82uzB8bXP0xSQY1iITtCL5rI1rIFu
d+yhI74EbTEvxAKx3nDJ3ZSdtwjmFJfR+Yl7K7tpN/hKMffA8lBWPTQUkUGUgU5e
wG5RSKNvfjWs+tovH5rhlScFkRRt7pcLwoOgxaOOt+H7KH8JptRVKs/XwwFddbyW
UNl0YOReI+sJ1agtB+ku3MZQcEd7hJvpfNN/PeP99tYmm0IY44vWvkK5Jd9u02RT
tnhexfMSTNiwtJCNH1+yxT0eCrgLAJzhAEMEl3+WhwF+YLC9qnB2xzooGIFnGLHn
mIpQG7JIK3VSqHy822RwEp6T+0eB47bfhsCbMwyToAZzpk/ss+OE/pDFRcxO9Pm3
z9K7CAFlQdzEOpUIHF7xOjeXqXWDD1FULMH3ktFLWsI3KThL4A4vszXMfIqWx8Km
NZI2ms/hpSpbUsSnrdtWVE5yq2UkM5MgH2wT1nFbj1NqLKIOQUdmK5eUALIYG97y
x1mtm7QcvFIJOu1HGNAcK4AHwm47udYyPRrBxv0Rs/e8He5Y9+PupF+nwEx9QBPZ
O1ayYMI/rtHa1XbWBMz41Va5YHH9MuSGhiWtFau+0VyM4t/jIpE7pn3bpYpKIphs
+0hXXli06SFX1rL7FEYqc0mqgLnW2JPMOijxmDROLknACl1BRowaAZD66RWezySP
3poa2arzmMpXo5AwJZNdoKichkJv8bx4xGdpGvPX4N8nG9vl2YnBsb4sEdECrBr1
eM/bBTuwzQWtOH7VIQctrb40eupRYIW3nKp4mGtXmPBn0kEBYXX6KMw3ap21+dEO
/FEFvOffU3ETDjSCNJzVjEspq/gnYxiQnEyxCus8WAMhCI0xneCRiY+Hq8JCQAR9
GmxnbFt3Biu5yWVCCUynlgdXKRjLFoYO1Dp2CtH96y73PNXQi9Gicn0K7gpQfBF5
mLhai54UwZPZgkgvTGibEiYDhY/40HIrC7JXq6RQu+liBGW0xrirnPLIghGa8dk+
j6SZUM4HA3apz590WRDZUMTxn3mCUr+qCQo3VhvpSxj226JHPMjnrPNDb8QGv8qu
y9X8MNUG8rEXn0A8An/SPzsEBUPIhUCPIh2pZUriPHKcYW1laAOxMetBOCj9nabQ
6uXe+jIjo5KakSD51kDp9Isk1Y7GEd+19Oiu5xJVCF8Mk8/5eZmvlRUxTjS4/Rkk
erffM/XhLEfp95k4Oye4CNgbtsVBi9K2FZheLJMNGQhphm3ayHiI5a7vPSUJi5Oj
m4NVFxqZ/XJGRLnc2iU9ZOOuS4de6cX1BOPBX2I4fNvwHKq37KhGDzKviJGTQWy+
6j3YAH0omIQnYw5HcNwblMHp+l7nApIZIZEvBqFPQvxXaxB2mIK97clEpUfHg8pr
6RQVhmuIHUO7n5hL8RgClC3CSyjdVR2wzP7LjRTxYg1PCRqgr0k7ztxeLxRQcc5r
bkI51cuTLuB3Fml9tp9LtqWcTuIAsPbE9qwGK30Xr+wDOttwaNT7d+ueH1J/cu9F
Qgnxp+7VTp/oCcW+ksH2efmFZ3n2TxPf8zFdnqFwPXbOy88qfcV/p9+JLghFEt76
dYPWea9AaJRSVxjgEOCWS1kmxWLEVA5HGznUF761uja3EMx36RRaJE9ti8EEgt5x
d1h7f723UNKQlZ9ZoRQtP6RCv4PtHikomTRKFriYBpf5le+4eYCsXls1GV7mTK25
ZnmPl09Wp4jUi3VJI0WbC2PKbJeV0EwSbpFQonUGfptJ5qMb837rLff6h3HUZUXn
kXmu/CV6oyG4+68zUVLaD+n/sk/pmZxCn96/sNS5p3o8ZXxSc/TXY+9GE0ug5rOV
+sU7vUFzZuIoixRieveXnL+GfB9ODCuvBolgWNuWjpIkwI4ryUo7NjKQ5s5CMTM5
Nqblb2vn7nsYXWT4zYlqWqYWotRTGS9ZV/NYe5uodmOsx+3dQOGREhmmL/nfSEmV
exDlbpq3wwaXUi6I2J94iUbFt92KTqw4le1nR834Iw/rgJ6h3ibnH5F0qjP/dIrX
i8374v39TcOciHkzwNs+7h8yjjdFs1pKQaQYhIJ7N+WD/+jp0TCh+Y4ENBjCiwEd
PH9zsCPlI1o7WUca1KzgWLl+oXttdjZ231JSZpBYPBd+Orzp+HI2cc27ax4ZfVrq
L1mUllU/lE9cvZU+x1G02EPVLx5IwwLnlBwmaLsgayfNvUG2SswCcj7k+VpCKx18
mUqakuBBZIbo2smWqOAp8Ag0goaqGIgYWspH56jVDOj31nIqQ0z+yesf/YdYBsbV
fM2KNiPmty6Fu9Ks6TQ6eWwMrste71nB5nKooGAN4tgVpzDPx4uhPTGLXVXCeDud
bgikg+eG+MgmAEZa39sOm4dpg4Dip1y3yrF3WWXPgRbk+r3zElIgjvR3UPoe+bnq
bXc+hYmGDbopfmpZCLp/uMD0FDxY1i6Uv6/7LUF3P9LJRqftM1H1O2siuP9wYE7+
KlRZ+Uzi66jhDgv/yVFddfHI7ZW+OjWOONStqA0nRpbGPJiiSpXenXUAQwvLfLXy
vWwcbTQA0pJmtuWFQpstwa5WLYHQZSClyk4qtvErRfmmTA0AfMHbTuvyfxk2ue8o
kT0Ebx61DKFjXDtNb6nJ3wfw9D+w9804WRxUGrMJOw896wQr2vU9xg3IDu+2rcXy
pfQb1ppvJ0XcV0ROaFk1k70ci9mYX3NPy/jAMG8NYzJ4NxX4dLK6dhsWm0tITqa0
M6YmG57KAQlkc1DfWWbuLB1++3bNyoQp/4q2MZXiad686fM/WCXejGDFFkMaFhw4
mu/1OJCNejB9dqii7tDk12jDc6ZQzs/2PIwZ+RPZWMj7HK4poAw2r8yjZsE3NW0U
yP2SrFl8h4+TXOKaT0ExbYQe9IFTL7w5yDELeREBHQwuU4qd6qS9ulVGyleERO3X
fZ9OfIjQCrJ7qp8gTWZ/Dv8dJa2erLpMUoa5UmExgAahoJuTXpStnendN5hhztxy
WUIGa9CarL6brV36sIrdCVI1+MiOqxXB8hksEk1f2I2SFiBw/rIggpk3PPoXosla
EbNWUreKglf/+K5eQNkyfUcvJJDw7C5t3IPKpoCqWrLqe1JHHQU/wKsMiNuTzZwa
OpId5VbcbkqtFn/44LcoT5BjCzocjDPeVXw2jdQ75wRvd67VoV4fACLBafPMzAps
33H8YUFmv0Y0gAaadqt1ekzu3/7ubl7L6JTC24vPNzG5EjVEJUQSoZJPDHCshPan
XWNyR/SjlglkMLt4sCzpm+1X55RHNNA2TUGGl/QzNo40xsqVBukS2MWSqb6YvNkS
n37PV8pn7vHVYo7hezcCgR/LnzhUZ7dvVQsYaH4xbqtaN2H7nZBVMYElmuw+3yME
fb5mcXlB2CubXcE7dH+kIqAmnOwH+crCepMmdlTP9pjRplG3OWVTsR3RwEH8bH3n
X4Hn1D79+tiveAa2fTBvoHNucTHRPSw80Ed3cIv6GoEZ9hd1U2RI6exF3nqLIuM8
XCrESIZqWhD/b7j6/vcDN1BH2esZeJa9Pe5+AXvlvKbJJY7OKRTnfdYlhRCEnPZb
uInJCIHt8DtTvGlHeZIkKPYJ//xvc652CkeSWcXPUfFAPX7A0SEHDfEzvC51tKJ3
ar2IyAJuY5Eeoe4Xt5IT49kUOBYw25jMTj7L+YMNwZIXLA3OaChDn1EkA/oK7OnV
rwa8BEfdHw6WvRkxx2YU5Mq68cyojHyXnt0O2JSYEqkFC2jvs2IlkL7Jts5MVv92
uBIPuiQo001mul+Pr/wNAZC8EX28fIrSidrNdaCGo5W6QdLjGwmKJyq9y9gwjFhj
BjULScsiHPmkZbFOil2vFDrI7v3KiS0xu2sZ/Q4ACm3Z3/nbV/Xg+OPEqMheMZYV
azSFXKkH2DDG23oRPQalwwpEuqmGaK3I1FklyoXLImGwPND6cv5Ton5NnptXpHBi
XFo55ZFevl0sJRg6FQ5xObEG0uRRAVRgztHAK1Y5mu6H9yR82yVK3/P9ivKAnZbM
2/CBMroKNP7SPdYyo7cAMBuIbaUSYLhJEc1MNXgtpGPmak1YFqxl03RAhMI9zyAV
I/+xzh/qlkUN+Dzg3sRQUvOsp3DNlMX/X+ks0EUmMTPZi0r52MSzVf6bjF2/yx/G
imXF6u9pPL7hlroE5lARhLa637KUQo6KnZfqxXowViy+N+qyAagVqODDaltr8wf6
D9VXjxyA+xvs+iiK7Uojv41drL69Kt/wVrJezGy+Ft9/kOBE5yD2QP8VsP+ir5Mw
eN8VVYtHzZT8B1ywt+iLPkwDHOJw53T5kVW4BNuqBwMoh2l0zHvFe68LDOxQDou6
zxYkiPrhPKOFRZYRKr3GPxR/OahEkvoXp3jWKei2Lf7+uxQrM+oiOcQ2mHo+66nq
wRSaxLQNx7T2YuBzTj9U34SDhlozESnGLaaR/2cnACNWnkaT+3BJvM+d18UjEFym
av8EnU31RSU6XfrdxUk/LXHSKD119RORoXLBkzvSCQK2cWN9Ossd5adNuqLQKCVA
3HORH8HpP+pcmMrmwj3y2b35HrN+Ltv9MWMtNcmIpsx2HYazmCyhhTQLfi4JaHru
uAc8ti+7/LbJzoQ5ltspYA9qFAJS64s7xCns3+5jdg8KNGihUI+Ca4+Zfa0D7w8e
WV3YVDk4nbEVYMs8U4J+mIJOR79CuL1rQBRykC1pdy+ZbMdzOWGdJddGdzyPulNB
+z5T6lTZmoqOZCI0zDu4wxVfmIoulK2vMMHFItdVRi9gZGR3vCTdIQyh0/Aa46JX
CW9CVqGo3f0dn8amiR9TfYBX0UITSuM6ZvgOUts4h83akhjI2SxXPrdrOqOjTHTD
1Qn+ITqRjLOr4WoBgemmT+sBuQhfwAxFajHeXj6sQ5ApZ8U+fmz7eZjAyJYhQxYo
YDYwPRXuNTEla5gLFhB+rEMrCAubUEyiVTVKSeycwP59Ja/v9+V1hSfU4b+IUsUI
Lg0UmktAXMyiN9qfNZRtl7y9r1qPvGdC/T0kHHaoRJc7LACiHwIHdw/oRNMJ5zT4
sm7X4xWX9PScJf7vrjwOk3ccR1Xs60LjEWRq53rcrmTqmxwrJgKV069Rd3Da3K3H
MCyufgLNxblnO9yNaTIE5NBAQoVaRJ11DYHlUikUAJ3JkhruVx1Db1edxrhLLDYd
JKeZCjaI63C4+b3hb6v7tGkeSSSweThi/lSh0dQ9Zr1l8JFqulmn5MjL1gjEahTn
D7nce9pDUl4UxhwdT83uZa6PN2dk/HPwM23XtZa1UQC81OsvgMunQPOhHu9UcVGv
5ErtWsyQ4T6h+CUr7lyvJloH+LqJCdhoH5BREK4Qkx155OCr8gxy6UHS7xJzheJP
lFcBU65jZ74PrT68c+XshSJQ7ertneUlqviECNWEuuOyh+gjUncoi0zOVUI0sKUt
J62vUi8nI9NaLLrdshYaUYQv6lRdHZJD/e3qgHynzm7ZyqLwjA2CD/QiBscHAd9/
bUEwsepz6eFGnmZDjdsjlqaoAEltXYpb4rv9HrSn55ihO4VIoD0nQ53UBjQXnqoN
0gmxVYBJ+6/pUyXQHzlGX7ut6l1NlaO0PzqE5AdqGSd4/D2mSQOTLBhgpQsk5vRK
kXx8clBup6ilG6ie+q5XHqxmVoxwJVHj1q8Zp+T/KV0rUbPhW9nZrrrQ9Hjgmx7Y
p2LImh3avV3nLToUbE52Wbt3ui5mWmzzTE7CaMi3JcfE58N5AxDwBbCyDgAGUR2Q
qCi1/mbStLXay8xALGqge7wp2fLjdZzS3Tdr+ifQRX96vdS42EghilbDGLW0/pKC
jpIduxana0ntckXb+qkj9kAOgLH16one/3/UcnPDPCiYMmzhnjC3sFIH/IpOaTrg
oOv8v2fJqWsmrp1B8v7mv6yvGvHcYXU5B/SCOsPJSbegwrVsejUC4eiHw17nzMox
t7srMMdQr00bfUI+H9KywvSjtHHU7sHt3FmMgjPhRpJ7CJFC8lzQDnUIwt0ZN6lj
awM0AX7A5lui3FcPnTNC1lAqDiXgzukEYf2NeLeYl6wxS+ZRWhEglh56ZFjzFFPx
caBAW2vlnv6W6IASCu0rwFzS04GfYpCixkWDmYb0cd9dgGS7ik62x07dBJu1wyPb
Hd/5vxSfF/ZUDZit5tSEjHX3XHZY9KjaYlZfp2EU2mrVSsxCcTEFaMVCy6Ap/Ba1
u2P/A8xiiTF+ZE4M0Na1s7mRyFNIfkUml6P+7fxgMOFKffgOMW0KxcH9/BnxpYng
JPpzMu+hmTPHmaGVZbftoF8D+0YkJ04Oj3DQV90dvtJT5HrZjdktRSTxcPfN5dAi
uqQapX53eMiGpJN+zd0qVzg62kipRYEOfvbizYIuA7K43upIL6HNw2ZGru8v0+tb
aF0e1PRoNSennDX7wYbEy8hedQQvF7F3/Rr3kekrCAR2Dgh6vJ3rcN1YUO2uiKP6
4h5qqG4QM+i7gotINCiEAvQBBOZbfTDtIILFyYCRFI1uFtDIDlEup8b3cuXSTtp2
mL3sZtKKq/NyoULC6WZkByLEsdttVDhw/4ZHsyQb0CXJQXJC5IZkFDcQ3OpH/CxW
qqwyYZg0DKUo2ON5cgOJHuA/v3kxr4Qj1GlqjLk7CmyfZto6tYW+CB314UGexVLX
xdSUPpaGHjdD7/WYcvmnPSVHOQm0B/MJEw6nsm13XsTXVp9MTMOBKK8KHbc0D4S9
ZkrTXrxkxOfz4csSQoAoqoe4dtoMbyvYbbFzJBlQMAl7t8ZOBY5l/1I4Vkr0qi1n
TPAXJRcV9rkM4Dyw68Hpy0JQb2QI1X+cK5MdzvTQwACSR3oTrOV8EXorU32nglUL
NsTx8o9W30XGgMalu/p/sa17OeL3Jj7DWO3CwfWwa0HWLsgs0b/OBqdZ/S6guN3l
kJH4FkQPJkD3LSJTJKT/XKdHD8Z/Zhzv/hqLnZ0b+0aA9cUY73otg4jgfnDSBbbe
lpkc+j7c/0ziTql0U8ffi421rj8PRKpt4vQlEutVkOjyxGHc+0KexsBzlf5KGfW/
p3s1yh9s6OKiwF2cu2KL6SDde87Wfza06YekF4xa2BwWzKro+MKrM0JEQVkp8k25
Xi52atxjcwT3sc8G5Qu6NfrPJarAxgz0ifm9EHYKqKis1gOXoBab2w6sreyIw14c
qKfs/gdTs017/ZhFml0cqi/XoVGjQgYVR5ZgA+Ab+e6ZSdZwS+iDwILolVniwM0l
DahyTylFFkkfhYzMaHF0qksEZUarJe7oT8RaSkZGyAI8LotsnbODcCQikyVA9gQM
cXYlQIUy1TXdU5zPagJBG9EdZYVQzYjCJzDTNIJWK0nmB4I/dDA5LuRO9YmM0TBX
eoSCM8GzulJMq7oqeR7yme/4+mdP4BEl6DOqQcXyVI5wjxbm8eHFO2NE1X27/Mqe
UEmKqn1oyQjtpEv13LhyxlIxxFHUqVp1zfe6NlsBF0zd/VcuzSfS3UdVY9Opxd+b
gulD6u9e2k2CEadR7TIHaHnkKj4LPNysXLAM+RNwPX7XrTKYHI/s0fo/ef+FAVUR
I16OufFegu5Y1Mlf6VHgxip1SIHbn5QFFmwAlki6t1oO3NZwPAB4GezH2ldZ0RYP
hLhEIoMRFMfM0ZLJ0fqcld5YsjcU5aUuppEn3C2/i0AangpOSTXxKNXjl1EnWKJq
+IIsAhefICwUZqnxwu4mJSQwKHIBHjsj3cU7Bwd+TE0KXcaUNb7HxirPlBa5mdQy
ZlxF78fyrXRs8GSmxcDwkK94aZEuKvNZx/KF2M4XTGa/sjigT8jRESTX2aFDyicI
+5SfFQ4M3hadpuKIc93By30/HkZRXTbiex5rodiJmQ1yDWAXhTc6XJylrcCY64Zc
OTBJvBl76FNludZLI3e/+VSp1B3ntr1ARtuq1vdQ0zOcsiEcArNf9DYGxxzOD2aN
05yVcfuM0g6V5hTRFrCXRUDSvl9pwsXydRCZ7PL3spLxukrUdaUwleQcuRswRTl4
K+wB2ZyBWcXq2+g17PZecw9e67oE3GWVlcZAlLma5BXbdnc/UvjTdMFPc3+sslnK
9pSGu7CYArDxqzOmNdVWschxQRn4CPIQsPeyjHKcPHUPF2TCIUkjcNm1scWQBHIY
0N+caIj/LB366Bm/axKXG+geFGobcnMDAu7YRGbh7MgXj5DzkwgWeHpT3wzPF1wL
QdbmVRz0XX0r09iX6KVfSEsqHDhNkFRLuQiyP3qP+X/N/zn9hTR3JCAiR2R9CYib
EjXz+sCB0pYVH8L0qWkyosdJ/RSb2GhZxn36AyQlHbnxZyaLpw6H2+qI079YHCqa
cZWhcvURL0r81UGFzZkOplDnfkP9+dD0yB8IDS6pb5TGtls2FFErmhH04MGaEstU
qhKHA8ispdOv4gRysuQwIpAFkpM4PbveiW6QGx0Wg3nkRK46vU78Ez5p3lMR15cE
jQPs+8fCJyM3R+T/ltcQb8ueTcG/UjUcwRkxWaWZyv4yFB6/glkhAMkh+ZrWyx2U
iVBpNjrbXrZYjtqgVbu8uIUXqn2rV81lHXIYc51sXA6mWFwEWiehMxHp7hkvzp0f
wzM1Arc0J8OCdqQQ/l++gfVC89Kp6q7TgcI8jMTrbmeO7doEbxPpAiNdLXyPzq0J
TxeGDsJuz4yvLLGRSdKEBp0y8Ux1FhVRH9M50MhwEUIQ6/jlLY4uAaQUY44RoQpc
M7TErpO7Ka2pHWUwqeO3K4VFdq3q+KPhzw/jGAi245rv1er4HXUjmQjWBFKM1QFE
LjXfUBI7lonuPV6UWiwqRzhade0fRE63K259j10u2e/6FH7hjd11IU315TE9OHE8
ilIKW+zF/e73CYazac0ogsajfg29PlCo0Az5ZpnKbiDnyH6QUGSRkC2VPi+nB3hX
hC/8jA2p0ISe3bNaT2uEaczUvrsmeXIxiOVfz2IEALV28D9pGnxk65+ZCuG88qEB
1bnYiBGypuNPvnMsaSsycKwGHOt6Xcxml0ABRO7F1T16JCnJnFVvbtKufy5SunFZ
MUNNxBJEG9XqySi2CZEwhU5QHZcLAtBbDfLTJvviqSUuH8+yUORy3PaudUftgTxx
Af534dziD7IupEy+AETuZE/Mk9/6JDVoxWPJHKrygR7rwItquORMvo+xmPrvsi8A
fc/dd1KIxX1mknL1SLqqrdz2Wt4EbJS5ZLdZMJrKyZWvpUR3lfadVN8uXtyooEPG
qLd2mrfajLRinPowJd/iL//zPWlC1+thRvZ5hQilEHaorg3PPcWNUaXdpfDFEfPH
hIH8iJx92KqRvcOWNLcYU/yUMc+m776mDvbGyl4VkYT1VrMulABEaqaBW+cuFkZe
dQHRsroICuyVs+gbRdBHZuR0qGjBNEhQDUr3PfaOPg6IwOEXcm3ROzMGAQETIPuC
KsWb3NASdZ5CXxTSrERlgwJHlvVVVAaAfTprItyCB7xxr+bg99X6YqMRaIiVxaNm
1BZhm96QWdVzxKRWCMD5FDT81b7XnckK8McRXh3EZXRHmrHZrB8T87MM7vZrbp+e
Pe4WWOcbxVXfqRf6p2Sg9/bOFAICsaD+2bZF9zDKB59FAWCvVkDAXNoGCxe41j9X
RgllbNFo4GAYWm5PmjASo08IezWTiXMK8Yk4UMnHQj/PI50wjxLuzr9apJ77F0/p
lwifw5mkHa6KOjPmG2BAdve2zMmxop/Wj8G31759FQePUNXgBtrw5EwGBL0lG4AN
KatwJc+0t5bo8cqhsoY7wWKyZgTQA5Lfn8o3h+pDIq84BFxRDy0I07Xrx+Z8X1Cm
zXXu4WfVdvgvYw8xkVnyFLKCb+1vi/Gmi9/PzPZQ20O7l1Vs+UNkbS8ncP9ooGhN
orUenM0moZ2sctdVJK1e3A4zZZ/4kmEHCdmecB2GK+TH2WEJA7j8Ys0uT+Vs2aTx
5fLcW+xbjd4laLQUm2J71m78Qj0l4Ivts0eCzj4wWiD7vIVPHB4aWTmvPZuk6ADL
Gw85+Nnl/BvsfcNj8Hm3/0lpUWE46Ur1MX0fAdBnVbj1UAfKsJwcmby8qNlR9i8F
HzvEuXE4p4PKPBMAx9slYF64eeqOvnJmIQfnsXrLM43E3Nl9cC1eOKO+KnaWvN+B
dL1SKKpjiJsjWbsO8IwQ1gfiUZho0TVpBW9XDtYp3ed6mQZZlEFGyofeD3UWPvPX
oWIDxqhVOp1abCaw0D+gheCGhCRGYUbWLkV9OoIB7eQBBt5JzzMqGFR8bPRN0Dy9
/OZ4c6VqNfwVrcd9a95EgpelESRSkytr838vpXVfe3VVMiI8Co+pzXllpdVdM5xa
EHYdkVjRpn5m2Ghi+e4uhwJ5lXMEnaaFUPx7lE12bjHYqzRk9lt/7yrB/JYoGPuk
Lgl6rzx/XTJh1Bcnx8BH5PD7wmXZCoMfn8Up7NH/gdBYtNfQd3q6SuvnbcdIlLa7
GE/rU2xmFXWJQiLC/KkZXe+MKOP6HBbOuajWytl58PFLR5hwhFlyAVFO7ANaIzMU
nE8Tl15X35PwTjhKjxc2bbAEUutTscBOopXQzFpXRK8M2s68hR1hxoGlS1pumaW+
/PePz5H1ZOmCiuykWEkBjvhmtOoSEjKMh78iLEi9wVULS+22jVPjRDZQrKiBngiR
bU9lf4uFqMS1VGEAPu7ylodYI9Dgwu+i2SCelRn0pYbyWJRJ/qKCWoERBz20pE5M
CyWanD+9aBo/QcSbiswlVDwVjuU6YWEt06oJ92mFVLAcc1vwog1fILYtyd+eYDd0
lswwvfBfz5r1b/+QqB3h3Rb9xK3afHvjW6kHJMMK6KMsagd2yFQiTmvxhVsIpiyP
eRl0POmQb6eNVn9wgSl8pCaMlmYT87eav7HaScEfXryYKSD5jV7Qw1Lf6aXpHLL8
vxPv+baTXK9U9tu8wyYJE1qsJxblKIe/zX7EIy4+/bWxKmGjTxLTjyFd7tJPoVn4
9myzqM8kVjJxscFK7SQMi84Xhl0PdO4j3G8cV0bqwiqT5m9I64441m5X0O81Pn2t
3ghNemN6qWRpG9msRXMBl/bDx5T+qSsjqz0b/L92Szfs++ZcBZM6UBJMCmkyDj7T
qasbI1HNGipRdd2T62ObnPWlnumydNAeSjFMfIzC1poNqFa0A3AaaV75DVIX+JyD
c45gwxNZ4nhbTmfq3VK01ctU2/OH2ZLbp6ERaKuVuCOLCDqhSn/NW4fk/uLM2bKC
beGmo+ay5wk+q4cf82wa0pyjY7e/N3kCPhfLk0o1W/Bq3FCEF1p6ITdsTtflr1NQ
lCco9VigYr3YHvnP+eJVy8pOamF4Zij+8b51AoX+l0tKNRT9hHUIW2aPVjveTfTu
eD+Wr+BfoUODLcGjI281L0bkcc4PPb8guTnjK01UqBefgMSWcxVYeu5L1tF0YvCs
5V2OIVy2WaI2hdyvnDutfyWSmEurP0RpibdgPcxzmtXKWeBpi5Zj4KKyL56uQpjo
UvrBGUMpV4CQHytUSRjmL8TRbRkahmozDGr+MJ5TWPGihxMrjuh0lZe2TN8FgQxu
cbIWtLJPtTMQ+kXWJCWcLUZvagyScFTidobgGn8pFJaLOYTSXPyohEg2afJNOSWV
eds6KOH7M8+aUbnlX6zs8KgHWwVSg2kewUElEviJX8WHlUvdGgdaSzm/ISX5x+RT
DFEzRRz21+KjtjfwlCajjHBmeITvk72pBkb8LalVXFK5OTmOzoNu9svfZ5g0XdrB
o0/DVKMpnv/uRy/wRtYCLRgt9V8FUn6An+liy5DX0U6K8wt+iG5Pi18+he499v9x
Ab9J4UP/l+lfvH6hnrtw169AQNcijiLtA1caXSIkAn+Drr4Qe7OPonkQggC/gfx2
Ad1fLIUdXgO/vIuBn2OYZveDk/kyLtfFJx6wAphnWfzn+6SaiNcOAeQUAuNgMwcr
94t6batQ022Lc6BxVVqBW7fMAYyjlZds1GU7fPjeimKTubBGKhkYPxumckSCi+SD
jYrRybjp4RxQ6Iji9HadEuSGJAQh9eH5h93B8by7h15agC3Jhg6phRG+6SmTmBAX
ClqHTgJ2XsbzHRSuBAm63Oo6LBoECkzmFMdQL7YJc9cDI6tZLG12ZQpKhI84LPQo
ed2MkCSRdJEPlM72sm1coli0kZ70/4mlniixW66m1iET8zNksyLiEJNzL88+BZkt
NFjGHKoIQOzxZoqzNru29NUdPMM+1YY16riBhCg9PgYA/5nSoNYBbEgV3xQxMhDw
1eNWBeWoJnvR8FKiwthmkrndIyUO3clzFSUSLF0TAV6FwYlwcKXifZbqawozdJr7
rSo2oBga8ETTyA0o06Za0dbKYECFVKKwuIR1m1ygrvdnPsZ6jkQwd0Gp2t34Jt+/
AT1PNEppxniYArafMoLTqaoaCMhQ/6NUMXtQFd0jtJYJiP5fOMzDkCoLMY5Vo+8j
Fv9wERxTwSLpEgrHwNoJM9X/2W1qKT2hu0mAWifJVUkVvbaWPkdFTiBzVNnLiO3T
P3+nyx6NbBYDUTi6jN1KEsOWEyGYKURcHzUCSkpXLIWMAQVsUGfhQCYsqjj5WwL/
cBh7THN5jM3KBPeb76LwRohIiirjV9qq0fz4wZeRvhv28f1yMEMvCSF7fYZfjFKt
OTzCyMF+eDHyUwt2DzePPXLAwOuZbuxHPjJNIozP4Ma1BPwfFVrqjd1REmiRJywg
JBNK12HZkesSV5iG0OwAHsMtuyedqHIxZ5sMKuPrtIw8ABiL9yrxQhxoWIISYQcS
tfjAj1Hib8HoEFlfF4dh4LK6Zv3Vj1P9nad9mZtHZgZ6GXrakiOBgI4PsIwgtPHu
AXqTi7U2j9q+cR8MrELxZH/6Q6GdVRjhrLbeofKrGQPWV7mvR0YNSmHfQVolwgrn
Dxry6kHSSeYrE5KF6DeF38fNU70FwFCnApbtyof1qJW7CVMnvxvegd87Fyck0W/p
5c7KFcqNdIqK5DctdXVTFbtAj7ctCmrbYcGB2A04vxFygM/iuIS5zrFE9f3DH+va
1Yj2HPzYc0+JCZVWeYsptIPpeC1OOTcwkh09OSq3UFRdKsc5TxML79kT2n8z5hSM
Zc3jPAuyYZB7xvPFRSiHYJ5O559XCItFth6sd/RC+CYbx0KXfrDkbd4PiTEjsSY2
tTOC8/mJ7E6vBJf7S23L83hYwvalj/tva1C3N+D8ScrMW1piDaTFoEb91EOrFrCW
9JyBZ+Q84ly85o7Lj/jeYQ0OG4aArByRX7WD1Vy3eDGTk7oguK3Kx/noOsh09K/r
0uEoueZgVnIbZ0W5khrbTL/LgkaIv2a0CByDapOiWIpv0qXeRWAUcSFJdouMtGj4
sTmaGRQuKan3sKOnV5IaGuBSN/D25NZT7n83pqArvSyQCOLA2v7JiF6AZnjMZqvL
VTZrxJtlATHlug9V2IXaSuiNCqYZ316osaIiDxojyhqdo+y9MmWfd5j8KHL/1Tbr
8zLcZ038juWf2oEGtzNrRto4F30q7AIf1+DTr1UFq0fDr1fzpgaeBIDV/ChTzISz
kjq1X9njmr9kw9b1XlPjqvgin0wBvkP6MYvFklgeQiDoG96B9CxIAb1p7BFqbCfU
W659HB6gT6K5BKcUxVbYGhGmqVvqfaPzFEiirs08w92MDEEZlVkNyaNeP6rAAeZS
JotM5pb6DAi7XYeu0daPINQ9szeRkHLnc2BJaqmBowCn/Bu1thUixcM61Rouovsz
f6kdXnZ/uAn5SHm685eZmk9oRb7s1pRP5MqPlw0PEyLidK/lmvxrCH8gpHX+9NyV
tlsrFP/X2IVFkfCYlnncrBk+B2ilsw5l2EnY0uKlOOz5D94YCJ0Gdw3BY8Ptbj+K
CLpUd+pQS1zCTPg46oLS0WrpnsqpOMCamqSpuI1wUDHpU+jPn0dd0pMfPFOa6vZF
ol8tPVFa89rhj2pVC18dvXJyZZ7jkTKChFV1KtElav7+FrDWtBkPp6lzskTiiZE/
hRDNaTuEwfDQjBlkHPRDEaVvMOT+fReZQNkAQU0jSCHfmzzmw4hsvLUk3xcnVJqB
XmDXGTJFxtNWfXvnQSVxcOsmZ/C2eliZyr8vtmzg2RB48Q5oj0blg5pJ8Z39f26/
8THj7jf5dH9Ey4kMZHfoFEDn5YGPRRZcXOnFiGv+GpfLnv0JiqcM/nLP4N0i9UiW
7qVCm6gkD+OexztMDAgFPxLqXiaAUUHTTkbxHJ6L0VBJEbm1coa4WtBZltu/3Zxn
fTnMqSRuSXeBukw045d4I0CBQHE7MEiOENjivjVrZmHYxyfm8b2JmweODsGWdMbq
a9iWz8ijT6zyAu8BHYwiCj32pS2lCw/cble+i7XwuWSozyQv3u2ncIuvJ2izhdxP
N5Lrjx7srkj00x5+WJcQN9uRoCJf7NZwipu1UtHMlclGpOjPMCkLbdNrYG+7xIB4
vhhcxLKoumPV6NuDSKbAYYd4yO35H0KJE0T19V5zTadXR9e0hRBn/GyI6XS2NogE
SSIQNdWHzEkorjLHQQ2m1gMMli9rQpDeCOP8xfv+HtOkt3x4+Fx45DkyS4btIOTd
1wGdcMfbzLIO5XVxxgDtBMONz83Ig+W+siynDqrEhaT9+2RSSSEsFahBGhVILQl0
2h9/lWRTHxVqrM9fHWVTFfmgNaqPYBkAPdhEAV9y9hFe/OLrPCr2ZehUPdyKoQ0N
OrQZcNWvMUxeTuwfkBHkWI2cay/MYiCXWaoy3fg1srPA4psGqfKDp3luqiXNkmui
LVgCnCC8rrWoKW2r3cyt2s/Slqpx2abTtkd5dDoZd48+rtMZ9V6uFvb0yVIvtz+6
4Am4gsTiGZP4lSwOSpBIQBPR7FuS4R71BjK3xRdcT23+KWWPvZwT3f2HntGnWDfj
ZOuM5l/Qp586i3T87EkbVQ1X6I1jRKP3/4/MDBhrkBXcUdeE2eQGTg+naWknmkaQ
Ns3/6TsgB75JdRmodZnpvv5oCt+VhCK4CwMoJs1Rq9C1Zx87dXuoKLf666bqj6k4
rYr70E1if8fiybWQMyfDrUeNHU+bsZZTfWMzjq8bpizTf4AFK6WZLTQvYX+jtwi9
D4rOz09wmF3dYgPztJiOM1mLyKNXaCNQCzQiCe0mH7auKzkgAGGAYAkxnXrd4HQu
4Q/VZMnuUU4nIZl818WZtb1zFiJ4naGMUmjyLFyshfGKkOEa7h4NaQwEcr0Al/JG
tRXWjK421b//PILBqkaMf53yjktl05X1bl0eMWI0SjokDXYweKgCcyjzZbDrvQCM
9Y+7ZWyf9Ec0VSXEyOJW6dzgGR2NFiX/o96c76EKsQF1KBZ2ZkebC6XT1U43Ooph
Da1Kc7J1SnQyKlTN4O6rLwFsXRcIsCZgVgAZ6VRB3j1lhj0EhBjNQkfCH8VbdWD3
dvc/ZsyqZVh5sw2axJhjOsW5163IE3yHwufJ+mAw/eRKncPcdhQtIVO2HobBpx17
qIpInJzpJglFWnL6g5PSl28ltYCUfKasYtFAHDjmhy+/EbqDIhFNwjxn8U8p/u6x
T/jA8ZMz1KZ+qpp0rFqYaESiUtNIVei9f1QJXBnUNGlKu3JpeXILsUNoYRkI7f62
0TbWX5D9YWIQiGgn1X4OKhkOk6Wk2QskZZc0HpiOOciIW7fY6YNXFHpcNustJuuv
gl7wi+ybWKWipo1N1FoVBbmQf4Gs8EBBYR2IsBs6js8MAzQ448pIvwmAc260PLzk
dsJS2JfHMLbu00Mfz6as2DnzZIg1m6my7VIqoKwj1ydDLBYm5S5JVibs4ITVAJES
YMj8CpBfgHSmZjd3nbyRhEu2l/cTDqONZnSHg5N1mcG2xovv3MqThtdAfObUPjqK
zoSixOZU+SeovSBxRuFqDcC0PMs05qxi3xbHET0XN7HRfZSyPVfkTpC+CRZ+rbz7
a2gg4i3g+L9AkllF31OrwHGzrpgzl1I+OkB+92awI7ex2YZ2RHK+1iGdVGXPWU27
qIwDJRh+nIrIvctaDtZPIV6xxIGfCthkcAxMxbJ0E23iWJSU7tAgwt73BomYtXft
Jq4m+DcF8aWE82op+nZUn3wLAi9VCuiCErncepAojA219fyyNPTzgunyX1xkAGCx
17gaFqqNVat372Y0L4cclPvnPZrTlTMiRh4bDRCNfRsEiBtEq/BVkGJRgZmFbksl
ryWf7/fr5WmaaxzS/tsF429IUXJcYTjhhW48raw6IZg6ajy3ADN4BkvNQ2i3LO6p
i9qkoXHVy8q7jnmxk1AgQw73jo0j+eNQhQiZsxCNfa/AVBg7i5HDaZYHBbD1e/wG
M8AmdAGWZ88Mu81EBAeoIiIDbqXBi9sJvlHpjpvZndUkqbzpqfq5ZLnC1AxeN8+k
085BVopKZsC+kMzgWIam6kuZOjnEyOcqGJttUw8zqIUNKfdlewOCivIuAD34Jehh
Vq0fW6RR85ofHROYRYv89zohaMBX5X1LZMdJRi22gs+vZxSJKWI1enzyaP5Mfqeb
b0CUHWKnDFKJaB4qmQHSNp0eDEYggKeu1V4CyhViJWrwoHXTEjoYPGv/LErQ0wDk
tL7AVVtsQzUzVMYfXzPOmUud93iZSYeauhsAoBbooE33iN5NHP+Wj6w0aiUTRHzN
AY8ipV2xG5Ig28zZWgnf+kuK6SHNl/VGLgh45XDub0f8lIfmqOd9P7CrEf5jkk6K
88uiRP41Kg+18hnxs+z8IHeuO9qn15PBrTIqnKfx96Lx7Pf6Ob2n8JcjXwk3SQov
905YWgCfV+1iI7lzbchYLDO+8L/bHAmtrse7Oj7V+E3i+cvTgUyHRMCrxtrHud36
o4g3Gs3ZZX9KXpos2NT75nPDX20STsrm/ncpo5nUOibrEzUAhr8O1buEGO/361zw
kNCeJMs7CC8OCMCn6D6rT10ZeGx8sMa/l/mS9aMltO9c3buNkZak8ob3pDS3mCOE
Whf7ZKEHzlg5zXILE0phaIOhTJUGzVishZ+yNJxbzPX1nnRJgiWmPqACwREBoY/S
YIbEBcpO57e3TigzqsIrdnDT7lWJTaUSr/4CSMCCECrgVovfuQct3B/xYWK4tMTt
IFj2pmAO0E4Lmdtl7r/FLwNiSgzlrP4EHzwg/LE50rDoZV+/sIsPyEkNYm6X9qW8
tM7+YJNl/8Y22U/EZqWsZcoupYZrgHzRDxqos7hn2Q5pcAVsDMNByWpjfKpK8wSe
FcKykAOqOoPgLmcRE9gnMbJZjVUsFYii1t3u5kNOaUc1ikE1+mnwk4v8gnZAPQ7p
nse2+wqFJYu0bGjqU7SdlTn3IX29QWW8uRVc8DAUupRFgoBd2IBHZx2jkwLSa9k8
sEoH+5PBbDhdYG2BjQnlkAezIbxWXVXS0y1LY4/eaqD0aJ6lJsaa833zh0h60ErH
n/rA6kcF07Kj2ozbQVw3KRNT54Poc3opbBgFA2t6t+u6Yf9Bo2tPdGryTVC1qAlp
uHE/gsylvXmLOcEu1l9uZug+AmtOVAaXR3wD66yWZ6m11n8UO09pb3jOb6jVot7c
dZcdwbbJwaxz2EbQxPxW4nU1qc8hgczhBJ+TdF63Llg5NGK8OHs6qjLalfa9OOOw
AGeVNwzUNTMUy4mf3tzexC4UpaWXlgm3O8Tt/kivCU2bD7I9LWMpXvqEAaWh+Sb6
gmVABih5eGoxAg30WShmXjCb8u0k/hJfS5dRTrm3aJX7EEWEi4By8hNu+eStrK8A
F+YewBkZIwTybwi+Yx1MNgDf8lCjCmiMDjwH42znqava6bweMf9jzBN5OHfp//H+
eoUblhqgBjnVDlhY+zR2GGqJhNUDGmc5q3+aTHO/t+lwkUqTbcnGJFKaMASgq7Fk
+wQ03u8qMU4tgDsgAc1lxGZniPVg672JsijgYFZicJny+qwnjoMMRJO1Rmw/nLJG
Fepl/018QiCVOxa4q8KoQD/iegt2fHYyAOYJamNRbj6WSI22pwYKmK0xua9BbYQA
DQAF8nQPdf40KBmnU3K/kf778nMtkjkKjMxwKHiQq1XHnIN25a2DAqkQXxpSbOvs
rYpTIVlw2j0PXfmJ6FkpYE8l+uYoOLkYpmHLCPSXVo+mq/bIH1E32alZugFKd+3I
2S988hjc0sAWwVvTPCiHlIfkFw+qZvrMbwfIkDxtNOE631yx2PdK6DjvQUtmfOE4
dJH4JIxOtCCk5jhltm/eXWkD1P7U/qjn259FeUFQWqfRhrIH9Kvkl3zFoHuZxyiw
Kx62u4YRyJRtT9tlFcDNWjuOtIPAcRdaLzdEo4UXDOgliOVv4C60oGjdGz4VaKqo
SN/Gxo2KSBhFGqSQYhOkO2o+ylP5wHEOuGHiAp5gL0eCwOaqW/xeCppNNq3aajfQ
8XW0MKh8Vh1+7bmMS6sdRslGNymomzWCSw9XzBcBOgaoCS0eJu+9YSaKPq7d1q2d
ULKr3GHw1CRwugbfazlAulQS2KtxWmE5USyVfYCdETzuMtzToYkxihJKKBelN8Aq
OsVMLctwJ9Fs2rWMv8uuVKzCpQ8q/t81A3gq+hbm7WJcGVf1eCUpGQNiySmf8EOw
n0Sx8O//aqVRBBNE0bJLad8jCVnwtbJFrgpiOyKZw7iklsjcTlcBIugvit0gRYo9
uHx6lLc0H/jqQ3t+wUsuqWqjGw75M/ZeKQU82x4BuXcBbUTZq9aPc8pg86I9raWH
RBaw4HYSXTcaCQ2PMY1k+kn3xVo6jN8YNhZ3kIct/qikYtQS/vO+8j1OYRCW704L
/HpauNyRxbAHtC+t8yGDMlo70mHg/9roMDaaR0JmouhQuKMMtF3RhEwJUBl8y/jp
LaX3UArzDmhVlF8B5C9yQK+g3qye9qQLSNZQUHzCf/JIXbGuZDpc2+BiVD3vrrmR
XBGGbYoGNO2KVh30BBqy9Ldu5c9/epZl+4QR9+f5KBkfaxb2Ona3TH90l8BrpQJZ
8SZo75eFzwSF9epMu1jPLZTLkNU7uqt3Sa9bixblMdUqKXyJeKaY5oKtJtotFPt0
O5DoOdIvDk0I1ZZJ8fY1hsdcYymbBaRYx45ch5xw9bm5dXY9dDhZfBXaEVc2iJSD
/Z54MpJWeACVqJgjGrX/ncG7e6A/YK9ROEJ6NAFNsYlDMnYy0ADhPtBA/jguwydH
x4Pfw9GkmHr+SAkitfgXFd4V7RxHijT9D0x3IY7LOtbW/yXjCyVrfWl/yyeHncD/
+73nGj3Krri3MGpuZN4uy111YQHO8wjFHgGVaCvSic9SQrDIpay2y/LggIzegjZ2
Byo/UA7xGWCy/0G5cDTFK0Fu3Zh8RzVBcYy13Thrbqo/VuvYvElYT70bm7oiTGrU
WE0QcRBlwpA3Syyiat8MeuaP8up+xHl/7qFwJrZNA6vRVnWxfC/4goCjsNVUiwCl
lbzfeC3INOb5FI7ER9jc59wJ9UDobsCXbc4z98OmmWrBdA5Rt1MVQ2ikCa7O6WUl
LUdPnTnUukDV07ggX5JOkw/wLwQgezE1L057b4mTBeZyuNkzT0+hMqGkOWzp/+PE
4seoRu38cxwSQnvmIF75ed4r1aZL+AsPwb01iiFPJqCHaZIDFFOjj7vjlAkKhgUa
U90s3VGJlSOZK2nnCs/GfRQGQpNYhHWLwh6yzzxy6I2v+lDTyxEo3GB32cjFgAWP
BY+cmOpfHqLJanERbeU7j0bnVIxkOAlcMgnaXvRl9yBcOUFD9goZ1iK7UQzQiitP
t9KzFtHDi2hof8kw63dLdIvo8SDpEckSHIkNDa/BvN3W4BcGkjnZOWwezikULAFo
/Q9saQoCN37E7bWxD3DvASDKRZf7GvXWBao32fcnoZhfQMyr8Z53ccyIFrTglkAl
AIoF8Y1i7gKjRskrkfFok5wBSLOBONiAsxZx0YoMY8L+DCwMfysJxnTfQYRfQpSd
xfgi9bpfukwi8J1WSynOu5lYeNnmgk7cJCywdV0vorJ4XdUp5xpBBdgQ7TFHmY6s
wOtYyjrR8SOIHnSpR7mGWiS1eZuJ7xyQp2tFzkrpaPNJmUfptWwXkDUGMO28QAJ6
KLiMfCD8LmKZ8LdAKLuNfe097HC3xk/h02goh8hacZpo+oVHG1KcFo38FerLJsKR
m736N5t+oiMaGxVcCoyZIW3TlNM2O2yWdYDCXYHjDvlHDTwjFcqDTItoTC71AhvX
1q1CQM8OXPTRQaJDUZz/A1ni3KQN6+nZ/1cMeyul46RpofYHqMYfuf17HTpzuvX6
8LKGMjKvQJpTvL1Ck8CNdrfKpAN42h3lAYaMjcCURDaqPNOdMZDVqyYubPyr/BOa
qqfcAZjxcVttwf2oL3X5A0yy9GxWSWsABHQVxYTCK1SlBfK7IVg5w5FS6ZEYZQxh
eyDDxl+hBfJNataMixfh+/9xIpQxTj+VvmXA3L1LIYdOq0n7uezBkjmf5zVraB/M
nOqfykx2e85gkp+ANETqz4uPNMk4zeydypjEjFWM5pvVfaqMLnZryFKCfxAYOqKJ
7jFBImu9thheNNkvSA+ybQlsTZZY8gW3LhgnDQKudR/Y+4umncYH/qgfdbEEl+1/
pBHruA5xlrM0w9cbv0P25hIORZaTqO28cQn1pMrGARKGtgTdFPTfPgmkN8nG72DJ
JjJV09Acvrqj3qzMEzYNjM7MDBMamBTKBgfP/DkB35tcI3++hECC5hAMVJWTWtnf
H25/b8bUK09ucnBSH7/Jh0G6iAatvWqbQ/zUOd9ywCp/NlWBdGXpNxRUs+iXLfjr
JLG3/fjBI/2CSk0OdETR/J7951ZM3quBXwB3Eto82t/WhsWOTavHSGRBCpdan7lV
5xPBj97gYWm2Xnk/YTRZ7x+TaG9RQ+kNTxG8IXUpm5iudhqDzgUQse+hCc5KExDd
G4rqqseWjLIEaFKnlElq/TKuZmrBYcd7j3Q20nXiHrxNM9L6QnNEyMUn2Tki1dnV
136ocr5CZ18vKsX+Q3FQBfnBKHMupBhdzVpysFKDgJ8TKfAWUdUTKh7FAWpu3g1X
yz4q/h2ydb6JakLk5aWDMztsTPhPlVrBoVdYCcyRJjEi3lkGdATs0a9Uu26b0UEH
2nIWaBiuJsoyGVywMag1n4h7ZJ4HDtlO5QRy7uOOwO9cfxG+Q+ZRvh9CZYVtCaj0
awrdO5qMrq8XIXQRKyyjskBBnz2F+aDenIaNMewhjDNV7OojA92/DH9PYVu6Ld6S
j7zaJ7CTKlnnioEoUuupgtw9FmIS4tjoju/nG0QJOzu/EH/qckAyQlUfoQ2bsyd8
UbvmZbcEMwuiJN5r26COupKz3mqasAk0e0dQYib2HQPwhXfjjRmV6+rPBIHZM8xp
FgA2WOAnIKlM+EbzAPff5cGrniMzO0jowr5di3O1R9NaCcLiHSxH+yZHBahpLXvR
DzxmLOYjS+znLy5MSep8PHl0eGxgxu/4iZYKB7wT9EyTJNMkMT4wwCcombpy93Mx
itnnJPfM6xGI+hc1E3Z2g4Efokr+s9NJ6N/oO+HzPJMNRXx9cVtCM6F4rd7VfSlm
vUq1vTUyA34kmgeLe3xiTnthjpi6qke+vTz8F62v2v/F1glcenfoQw7t05A4aWV+
IyHkRTX9UQawoLujGSnG1lhku/x/ugvdQcBRntRToaFJsI6YpCSskU0DvG5BYxoJ
ieBPmuYZRVKRUbF7AIOlpqeapHg8BUVp6sLDfhTa0wu7whbN8Js73Uu5FS2c8jD0
fSVd8Ti6cpA8K2LtQqIr5Vz9J91BvU4rKavpH58laad0+a/ESmsSyVCYysDoXgaw
LiD3f5ygBNEgYFuU7Hy5UcLz+SDWwE2w2u4MLEQNOMGNXlVUCTPIUxn41nI1ee90
g7uRdbrn81FwPBBKEDUwDntQk4ITGr6sGOmmlI+MykgIdlGvw9K0NjXJ7PKlOTQR
NUP4VPk9ZUc7OSi0gkIXz+qdYhfDvKI9ILZpNcbW4Fqa0suuv+FewYJgRyjfOXP6
IRVbVwSQwsfYonn3WnfSRTYSCCZzZIqF2wt/4G1KfoNZRvrhK8czvjEIPW4V7d9d
M72rK/4w/d5g7ITiYXV+ivr+AqWkdGFKJNpCurSzxOvVJkQYL849GQCO3OG2dtcT
1I0zufMHXQ4LpuKjSXgwnyEBb0kaoBZ8cldyEl8wIRrzAxgi1ekk0I1N/T9XCaHt
PKlTAtyuclf2Pi+BhTXjHt7UNf0XHfHsHMvRomb/C2SJpuwzqF2OHLGoA+dHfdCC
dgvNE3x8M+uH28ggADJA/j3AVOq76cEYz73lQt8lKWo56RjrdZUv3oXiMDAL6r46
8KPh8MPSdv/84xcsutSa51mfnzpo+O5t5P0jwY6Qydyx+BLEmNgKQTkM1lqJnYKS
0wuqbW5MkPNzCK7Ii+USBH6dEDVBXJEZf4BLeDSJpTTU3evS70AmPqYGFxwgGwNt
TjalJsFWsZ3x5/vbAjidLPgS57U/PjAmi2042cD3H00e/DZyl/KAmCLrazdxJS9R
5IBTqZPULiY0EqB/OL4tnsDYUtL81ewr56lNzgZ2Sx607SmXZOJWGj3AywB904PV
BieZiZBPOtFOtZu+uxmYFGu5aNTDZe4hOykby01hvL/CFB0G9zrimzLcAO4ZqRjH
fDaDVfRw+At93Q1KvpEvUlsBs1sIxoSVVS5LTAOyuSSlOo0aVfOtLPqqxpE15MGs
Glw15fB74cvfeGtvtow5S+nJJL1M6vQjxB5b8ymVTeAHmhHN7FGpOd31ZW3yI3Te
uZE+c8F4dnavTs8EFyfE2egmChc+/9jETC+mz5Vkmwd9R7ADNfwP8FCz8MSJqi1p
w2BRrL+38MEPT6XODdm5tDi/j5tctVZZzlJ0UAZvwXnduwsRpKMQKQSEcE5NaHfT
gTdof84JqDXtV0bAfUCCgNR9HTEC+E2QgM0LQ9SylQjYtVswo6ebAaM+J8GQiT27
79S9z3syyPx/X51R4W7Hha4hhAbiUcd/9tRai/fM8/IwWYCSZuZV3dQQJwweF8f7
ViqNN3A3MZ0rRqM82qbW7cQsdC1ugcryVbaOskqXt4jvTBgjEIKNjx7SMzlLRy0w
OjKL6EH2W/EsPtGL94NYSo23YOneyC40Ysv8853KIXcvoq+q0Qrg6Pq2FUf8mFdh
q5McXEmNRmArxKD2C7O249sjaK2tkrkbbjoW6joat2jotwvzMdML5uNLVcxfeX7S
4hQ2nrPXyxKvIPN9S6NJiokq+lBtqQpqFmEoQZ4NYSUaLgn1gmGwiiTNWx1xoxpO
K5sQ6m9hjVgWI5n78ylhSLQA5m95s+w1LF178UOvHMNeTR+r6h557Rz7Wr/vvJgX
/xZGpmYnq45DTxnH7sNCNvRjfyurv0xotNLTxWeLvOUNIy9SvLJPrMqx02FOBkvW
ZAN9Ggz3SxxX00qjwkbUBUAzjAxVXNm6uFsrxn7fBa3yHgw41r3yI1V4qr11Jzhy
gNCQlCsSpULgY/axLrh06AuBY+EZt78XOHDHEUEJSKh8Z+YHx1teJZOEX/ZD1bXM
nz/eZAlCC9/M8JE91IRyPgluyD2GicxVmZe4xO4zdxxo+sV8shU7Yu/d/kQFz1zs
XqlZlNvYJZJj4Fxdp0zLZN6uRub977rhpC0EXbmwhbR50QS8a+AAP48R+bLXPc7P
54k5zp0Q6Un3cTInhYyJ9Huh9BoQRJ3kNCaw5ffunQnlVIFDP6WkC6iMwN/P7fAR
XF+n+LF/wbi7LKRUemgLJ/yYpmidp6KlNUB51A2OLoiVN5Oq9IpU2LLnHEwcRtM/
cPib3L7E/jRFOVbjeasEoEkNbZPb/j3MyjEhqlIHCXZpLtocphRVM+XT1ZARYrle
58/19WFNiJ+94X3GOpUsco6jzll1skwKrFTbcskTBHJ91blNf6zyjnqnSzLEljpo
BJNf43/suk63KESNcXsrEIzI3h4qoSFBZEBZImsUxotY2gFokkvvM/nKZUAa2tQn
ecYnGXtE/Ye8N6B7uVVMNgHa89xTzwFMAzI/8zNuJcer9tP1Y/VU4EA+DtOPjqxe
KTAugtjs3uzGUQxRi3cl61mvIrvM5qznsZTJungMNsBi6+UKHmSFrFyht1Lj9GCS
+33YZzmUFRX1VLxItjK1vjgpJXefIJB/qJ5Q4uRmSFtSGXF4NHaDKjvKnL3QPowj
MgTHagOr5215hwSVxRMlWq/EhQxPQryzpCoPnEWTtJ7w0J1sr+MXEAHjb0CagSsE
6lesPYOEZRnTq0yGVGTrGPOwwq6Cd3LVMemhq42vqH6AOV+AIXRbCHWqPEq8w9de
tydpNMXsOmpuy6DIIy8s2M0z56fPeC1xg4oyb2VUWF1Duywo/GYQh69KQw0/FlZz
qvxKNIBs4k/OUQoi+0hWBruoFoWhn7ZYchN7ZXGhoOZ5ySP+nhq6gK47exWAdRpo
Ee+44T2YPjkbV5OW6mW/mHMQoxbW1bt+rr/kjNC47QgCXbrWTOnSgrLcjQ4+kEh5
8VCcUZ+lOOWakfiy4r3xmH5IQ8RpjkSObuBQr0l+WLwlPFkS/b3oq1ojdsdttEqd
zX6r3xUHeRGbWCu+9ijW51jD50OS4+EZca4Cka9DyZSak54Qt8L6bb2dxj2z4URy
8+dpB8/SklQEX6qMH1h5JfNIeh8XgqI02FiB6D62TzgYmWO3hPQGkEUS+By4UVrA
kXLLdiZfYYamFCZGlpQXaCBJ4GsPFlSBMi0Mh/Fiv6NSjIcoSGWXGx7ZNgByAL79
RL5k+nQYYHZbAZ/Xmdj/8psPvyPgIybvMUwAk/iRTnOexs2EoBcRxCdDEFHr/ZmY
JCye+LiIl5s/nYVxARvLu5EKby9hPnF1PDkjuzsO/RYDuOz0uG2lgIH40BT0Rtji
ZL5rmRSTi0aSlXCtRxY+j+ELIY19FOrcdkXEIFkSVGVE0y2AiMBu3kjnL55Cpldy
tNZIIi1FJdFgNkwT/Wkl4qfyTRjFvLo4oKoFjf/cRAGqLiAvQHo149IR5c4frwGV
M8UkmNSsx3fg8CFbmM7jwwHB26imCbJ6AUhHJj0q/vM4fb4CcxAlZdTAnG5aJtJx
xvQE1uqHeErAIeB8zV5RFTGK6q2C8U/RHiqvAVUan00JKPWC3QOtsgLz7Ifr8/0A
Dj9iQo1UbKPZSoqKZKIA7D9giPh8x6G1UoYUl7E2rBU4RyTyK6lTSd9rybIeI6Ql
+pHDzxQxx48M4548YGcI0lQXFWKHb96cOFzoPdumc+Xh/YsQFUOeTSjQInZhgF+3
NqI5Amb0o98jQfvINIvOcCQh7/OCCor+PFC4ZUhnN/zs7XPtVgopAW5n6q+rRg0O
SPy6XQBiFJqYIbikkHiAV987Jlv43ao43x4+5p3vyjry8DTAl57fh2u0T1Eh/luh
uDLmNV+9f7ql+cbnrHqo+bE7fENqtT3DRGZ2fO/Nu7FHDurfiXGl+7hdlaXNaPs3
LZ7XP5PdbFrYfdAyElt/37tOxQ6FjeNxzfVMpC7XLWHJLec8g1DrIENSa8iBcUzi
bV4vcik/RODACf6kDCX12rsvEvP6dWsOyNpS2VKHEdshBUPNwY+gYqtTDxb4zTA8
8h3HeReBTxN0Kk5hB3uoIWrjwfoGbLYWBfeaf7zK5mkUtx7oWx3xzG7/UYQUotCe
pjx4ojKULHqq3EJlTt0trTW29P4pzulARIjdfMQ/XwUVyJGMhnRQN58A/jgcoKXZ
/bVP5QAqnVRXLQQIECVOyYWwkdec+XAO5uWi//JkgOWPMPdw0V2SYvgqj0PDV824
R4mDGD6LdhBwByhLIMTJVeL/fHd4nRO3Ytmp6bt+XgAVcZexdCgvy2ijjwK3lrBZ
+Z2FLs10tQLXgmENv1sYHCbWZJFj7YcLoseldQCwX0e17I7hk6mdKC/fMTH2AJwm
WamKii6BaMS7wPo5AgArU/Ew+OwlK5hoUx9sJfFpj1mv/XtxhruhFD1hQtpDYcVX
dU+meVM98XM0KliNoHdbZvGCDOWcoRDeEcplDubdYOWv6RVKGD2LH8gvGcX3pB6X
Dl1+78TnqZwD74etqHsa0aKikA+IY2sm6wFs11uPV0jm3sj70/QD/7zLg5ns8N2D
MY0DLwDZd/YFfo+xUWPny2vfOwHQ7nnj1QKbcBSCewBrI2NoIvfRuHMQiGnmgxS+
LORRhuGbGwaYjZnONdQApVpIWSfKP4OLCAwaUnajD7rPk7UokvqrAXnB/YutlqzG
2PqTV9PTD4P1HqVCj1mwRkuee5WcKjYN1dPVD3lgfS9dfztjMXA4+6P79NVNBCUx
+g2o7R5IFA6EGm5uI5yQ0dtKwa8IHfBqYBUjr0biMuVNJMJINknz5jwmr7OmDdWw
Fm7x57IYeR6nvkNph/BKZNis8NerPkCmBgupLowqWMNSL6MS1GpTsPs4zdWhIYOp
Yrok/qQ+EhfsoQ2MjKogELgXoy0tuZACJa8j6gwFuSMdzTKyxKcYeue+zDUfmmp2
zidMzNFGqGfZ9wHAb4j1I5zzhIW+0rHp8Zt3dXIZq52Ogrw6OK63SlHicIaDycOv
oKTVKfXdcPyZCwo+bC5ld+xFMARbtGBqsTVBTvKwKbNIrhTG/ReeWk0now5yYLjK
1pYznP4kLv0xxowdqfyAiEWnlsblcRb+E8gbw9f2dfEDQMDw8KCSw5e0j1Bhs7sx
1646m3g8UazramPlLnsS8pcGvId30M6WZyM4I5RwIWaE4sXT4q82DWv0E8OhYvAh
wuMl+2rVKcrNRXyOdwjo/1py+/fWR3cWX6Nx9iJbIpamxLElJcAHQYiw4Fuif65H
FirUPyAz0vvVJFcfyYPZtkBmivs9OR/sQzm77ccmb3sqKIJsrDm5QMco8f+oWzuW
e2SBU9LNakTujjYCMy+brptuZee8YLO11RmprCpczRZsYD/BMYeMoVG/ttP4+4gv
6BqQtTt6e14pDl5GOsU8hUN8Gzcly3l9UC/Rtb7lYs3ob/S7u15JBQChs7FWe/cu
syFRl4TT8Luo7wJvoGzDLCx98FFcVZgc3WE/c0Ap0U2W1mc5Ig++yKutgPAkXsmA
cbLPiDMbOXA730hxOGf5dpOV6tRWDz2boiHPw3LOlNUx3aL4wBcw5ea2zNF+Wqsj
RuRPrGShuVj/Yr+cp3yTtp/nm1VfNv5e3ZMCfnEpqM5zxXdbChZD3r9+Xc8bPB2+
y/HlGSQn+Pkpt8MX4WnJMus/kiXN1UkgTrgOFG/Q+vqcO88owsQsoFfBU0HeBc0c
PbxbCBP4wr4580zx4QsPdiRPCMb/Wwp1P2Jco/R6w6027pKIHbbVShBs+k0jxIaL
MkA+6m3B6fTMyO0hD+1nA+p9htwCBhad1zyQBQYOMGBVle8SrSzlnLKOTFZo4W7h
B+46VMt2fjyqKzU4onzsIVsjQskgWqNA4OPPDnP5bl3KUmfqDqzf0P/8Rgdj+3BH
vN1mWQpVsr18OpIVLZEv7Hg2u1N+FKLaWsioLqhBW0fm8Z3Ht3z403JI0jfOPBvP
a7N0DST6pkmk3CPUtSk5wyOGpN1dnOlOQk2QkgFx1xnl7yax1nwLvV87jbjLaY5E
HMZP41gLZHjSKslYzx/MkGg6Tf2SSf1A1dqz4Aq8yI4ouwBVgrZuYZW8JNms0Oci
oR8Q/LJ70tcx4nGNmgHWRhTEX7x+VnD/C/fWZeQrQzYiDJ66vIzhwnzwO8SwIAIr
Dwu5IgDpWCimc8/QRVCYe++3Zhgs/F8UNZ3I+ESe+Zdyl3+l849HBvdRCcQ4b1iT
3O4a1OmALZeGsu0M6wb/2nMDe1xsQ3ls9Z9gY+G0hzfSsnSls3bWI4gQJ1fMtg9Q
FnXvrIkSgQcfTI+hqYdzfEWXClKz3J+2gFgxHxAGXw1NqeqKtbGGcISYUJsfXS76
2DpeVAnlH/uC8FwhEawwIgHKrFvlNOvTdcximzmf82upG0OdLBM1IeOO7rwYjA4S
W99kC0w77PoE1qgPOEC8JwkyYfJhPlUBkdlYsFazXKH44i4DyXqxtlsBuzshg82W
oVKLy6hEuaBmIcgoST0fBC2IVTUqA0KRRKH1eXoApi6lE3HmKMM2wCoQMrWl+rqs
XOijWgT+pxSvLIK/CcLxiiBweyPuIVDIJdHm923zcY9N4M8h90GEN7AaWryQ422L
QDhK1QUyg0eR7A6RbPIi6mWw4cjQPs1+s6iVtmhcffJFw8Y7Z9jolmq8h7/TDlIh
YfQLtOQvm8jw4kiliJ9VRTvn6eWyaaEYjQNVgNRcXMfF5a0vStlJPIMegf7XuTBO
R+7iNE7i0oU00kL0Bxbn/1sWTfT5vm5w8HdXUBp2d06NvgCIsS0Dfy+FzQSXRvPD
h7K3IE3mKvTpdOcKiWYibrKpihuLMAe4nrdA6ROLuCD9JmcxTf7k1JN8ox4jua8m
dhY3gNdzJ73U3OCv8zDlQgnGMLZnsnxKdJDDqS/YbVA2n02T8NzFrQIAVYkl3NzQ
Al/UlTG0ADfrUQaJercYcXJxkh1TkVQhfKZLjo6z0jwyc4wj4DtGBdJaD75vio+u
ma3/pJrbuLjffSrhV1rs4CnGOd9L+sr1nWGYMfybC7IRj7CUVJ6TMZlWMD6OCtgE
ukqP5VfrGBAVrs8D/odzFYJHJwsHnFE5zctF/CmhdMb22gpKXso5YTF26DBon123
mp5wWTHXFbyMo5PzAwSCTP8KgAMHwQWtq2Am82qfTPjW5oltn7qZZ3lEMnvttl4F
N1xkiWVo8KcunhlkYYzQ3dQDjg5Lg77fPiHBzo7hb2hosgbEmTu8KHiKYlyz+nMi
Zef2I+gJSOKiMqDOy4n21W04i+yqrrY4W2HmSftT4f9/xayFLy18f76hHuBnRHIG
zHPpzX1TKnByVRkmzT36x/TRK/y5mfRIxa8rQ/me5sxnxw5q2jp4Z6TFhWJefJA5
QvrLpSSFyCNVPwge8SSxUKIyuPtCEDiUT8rbQEsljHzUjjOUYZn2yJAd9PcqF15z
zV9tDiu9laSXxd9/nlJ15YJdr4pj48pbWSNmgP9jd7MPJANiBKBE3LZOfyj5jNfX
cI/cMdG6ZeJGGSCD/vYpHr4HY4Y3Sr6W6DfyqM9vXEdGQnrzxSbNzKv8UcHBNzIw
X9ZW2sAupi55pwyy4nZ6f6cCWsHmlwayIlJi8FJlLllF+xyOuHHuzSd37cMzUKdn
ZRnpG5LUot/99l+AcOtacaSQKV7cr3Gr4c2EsNv0GeL7oIBs9Ys/uyd0Bx6SxRPG
FjI+YMj7uQIqxAQkB5ytclffpTpEnML8KCi1D/6y9X6Y+0flqPbnFirtmgVqTUjJ
AXS4uaNine6fa3rfdSmyZKQCMEVYO2FLeceNH6nualDHXHof4KjT6wZH8h9t75Ba
hG9Lfv/WBWsyO+T3+8dPFbHcOk+1r05mlYbzGuOgcpsMEP0Ajw+JyizuztHnB7Fh
PLEr8eMGocHcUfH7GV81ifu+EkjwktZWQNmnqylYfLvhOBEsP8qAl/BT+w6Rdd5I
BrLqvmHnsgaHk/rP9qqtfygoEX+W3gOmvocQsEIMnmU6DK8/Ui+xACcd5lak4MrR
oVbbcSlGZVZW3Y2wecoaPrvLfxS3rU6Nxu0o+8l0JZRwSeUkXf+S3YxUHtwL+e3Y
+f0lWOC0YYVnXn1cGsj+Rd39Xt4vkiOnWFGZeUY82pmGNxAl82D9eJHTYLj9JWUf
JlaPxhxsyT3iLoWYEpvCMJBk4BdeyUM9j4u4UQGR00BcfZVGuCI5EMs+otF0cq6U
vgYahhiuQeZHYPBM+IWPoGeMarEP6JJSCX4NElHkBoF0nuMOWGS/WiTvG6105h3i
PD7k6bLdw7uiKoTojQdHhzgLeQzf5d7GxsZ5enpIifZFuPGKncvueXUq/wA6WMzY
9T+jOyJjRQzQ5yF2NvnkU8VlbPymgs16eTcHgu2ecQaNBEZCT4d6lNaxjZMcg45C
2Gp9ZKfDg2LOh+vbkDh2+S3SDD/BgBQM4PaT9EYhQzLwxo5dfzWgmnBmDs2xNfhi
pR2OkM9N4dlmGSrSbIr8E6G5P2T9SyuYG52JkoYeb6wYbCQwuYQdqjHfQWH8xmAe
VzmTsyPoy2R7s60/H270sJ1W1RVg1RbxkQAfQ1CfsVb4OLO/K0z3nbq9yQ06eeaG
yRDtrnEAPAH8O82Hoh/wpFZpb/2eaqMHV6nO75dDl9Llw4GyldXvtNCRCKnpUBly
AslXmyPP0RQU9U6IgzOERf4l/rHf2eGb9Lhs6gQlkOKJDGLopbAKzb5D+YmrZcvL
koU8co1tMkQ6IyT7Lppj1psrH334Js1vT8aSi5/xD6tUexDMEQrQKzbOTG+qLyT7
zj2x31Jqf9UyYSP1nYfAp3YmOKLzXKY743SHusv+vSphfbyFjRf/n8IDrfJQAYAQ
JZSWpq6VJCUzokYFQpazj6tfIE7NuW7yNHhcuxP9efZYaRXBF7uVlQbu1ipAnlLG
b2b+cv0EUSCRZmh/H2rIimUETuvP3qV9nrI371Qcy+GzglyInO5oTEwHObp3rReg
tZvE1txZbOd3HMnsdhrt0OHPq7TbZJeIok+jndPhcCV2rULZXNL2a6iT+UnDr+Qa
siinU/eBfg2/XMHMEE2LBkgeIoOWNpmRELzUmkSMj9iaC+hx0Ut+0NSpmm6ysX4D
kfNB/bdSD4c4kDKJ0TcLp9W78QTM9vSVInd2p/IPb2SyeELAXpVvyb2duT/PtDjQ
omL8hRh7j2Ht0m3WHNdCHb43FW1E/2mLkg3MQ9Q2Krm/s7AFZQ41Xmpf0BTBd2Vr
bn2/gW3zkJnnaGG9qtVoP0TIUCjV8n2o2c3FTiYFI4xrLVzHlV4eZgraC7Dz1pAy
dg5ZWVbCCjhP6WYmthBB4sH3aBiGX/jqfCnjVyT021z6AcLdJeBr9YbEhRSN6I2Y
2nMJPavkYxVZ27K9x5l+95q7orZ7Omr8At+PJkixtZDK93I89kCOxGCjXNuOYT7J
i/oHFRx5PCbYeOAa4oC6bsN0fiGrPjNa7t4Dhf+UmdNl/JCigWqrDTmcYhy7Nh9w
MC9H74qdbM2/122JymJ0Ady1GPfGlGOgTU0aOgu/ceMv8BgoAoAOySi8riUisd3b
9UWTScziJqTZOdfAFKGcgwBlvdZhfYCW+sJWeeKz2UAKCZijwuhLM/UenrP/em7H
n3u6w9md3fktzO897H4+XkDG13atfoc2ID4Eq0inrqYrGSIlfMPGDdLHMny5J8yl
q2A7VK2iNzqHJf8dDRNP/mEeuwnlYNFTBIDCb71bLXCUkvTNxVrgsD5karWMthft
i22T7bfGbf8F0JXsyjso6yizcEfZPRaS0K6UFFClKmmxlnSAJQHPEHlN+fe2PyQC
wuP+IGGhz18zjFVrmAG0oiP8nS6zbeYfun8mQu6mLA+QNpOlJs26gzxRgvh01p9S
5ClZwNoa50WUeaE7Bg42+30QYNVnmwjNPnvwXsXZW1Oy9HDRoF7KQHXYhwDjqn2R
/MDC0Yzh/2NoelcSZ9e48b94fiz2CuGmPY+iFlwydH+bN8sZzsm2finwj9PcBjpz
6aU/chcbJ0SxYvHM/oge4YN3LoTebnjAmUwDRZYTwpdF7o51NJ+CZ1t8ajDCsJ2u
Ntd/khylz9rkumoi694oFVl8aZSufn7be3FrKuH5fLUkewf3d2y/Oj9zmEkAS/di
U9ufFkUpIqSu7eMeiKZvUNu9XgHJZxJUNX6cCk8FxngvSVIYdKPIphj2dPozxrzn
j1LZQV2CfzfZW7zDU1eY7yS0Yb9Rz2j+qYEp18XHDbr4aCe6M1qthLG+eVuP/sKj
RnXSLTDNyMd5ARWUPbrC6UVDjSgnVHNYiFPVX+tcS/J/Oui2KMMXKk3bYoegbFhz
GEbvMbM/EUmcNSu2U4KNX2ic9MhE3IKVUwptd8hn5eU3mOHi7qrW+sKU9hh88D7/
liMW8fiNxVWsuMG0mjHhN5dnmdXY2ctc6+I0VA6+lU72Q8zrEr5HeWc8J97oXHaG
5sZB/jaKLRWDzpF7gipLkR1ZO7kW/4GbXp+2hMvBtk9baeYaR0u1I9P2CsnEKxdR
cUlBcVtBGCFpguCegqWGYf/fu9ilXv3dMy2dcBx9BAyb21FDwW+KkIlrqqAb7sid
ZN15CWke6BVxzMjVYkmPMPayvBoKM/B1FIfwFWzh/NRgc6i5TpXdjkpNMXAYDYDT
yd5S32QFFi5BG0nkw5SSKg9nd5BrazG/aNHlV2iS/vP/Un6xwoZmg7SGMHhasBUB
HUlw+UYDVgwfBKCcQyrRA/qYDTG8URAxLib7KyRuIuy8YRunX5pFarueWdlj72V1
Wjfjxdz11bCiZbprKNeVr4fBdu9paleL7QE5ujzhNhrmQMLNcPyqjTMxHkNaeHhf
WG3PGF1p8k9OyygqBIkLP8J3PxY3cRm3SPfiSxMHnKMnTGbhIihkLIX11EA2t3fU
2ZLygHy4sKZBFpiYLDwkwPRwgpnW3caqtgwlntE491Kd3EPvdu234NYjgnj0zpD4
q5Tn0lJcQVrq8r/t3CxD7XR4ThCio9ti5DHpe3lYQTFQWBr8MDD1zvHifL6FYzHx
uyrwBKfArCBzArPIjT5a9z8iF7RwNa1RFqbZm/++51mOOiRT6Yo7SQcN3fesuJSw
fKRbY+r6SrloA2QinE2q5Awknw8bInmtb7G0XUDihk1Rq+SoKdqAjJHRc0HnOZF9
isy9znI8ubvEV8XvhdHJ6hgSYZfF0jtBRl/eyXBFwsZRcp/nrgRMw3kxt9zm1Y+U
fUP/HQNC7AvW6DCnhdG5QtvhUrwQ8Rp9vk5LD3RXbiq60Kzf1Ryj9PyhY95Axg2h
A2W8h9pghbh+9WTeBKfxJ64ZWTWrJdFN48lgFQ7TTD2KBd0CpUgEfHHDXjTNUK6/
E48dcXjfsq/dMgYJ5Wk7yDE5aJnJYq+XUkIKW7xb2Na6+rhtZAIygD2P/6TbsWLv
OKLMVK7K9c/geLDnTynDPaDkf5BKcREfMRLXho/kf5TJ8aoxvu87caaOBxeWMZrb
13oBCSkzjrNRviyGTciCjHeZWYFs+T1ZgtrMX5yjr+lbgkN36OtsyX3P00Yz3POH
MGSa/GbVVoZjOsgxp+67UkLdwOeuH9oZG+SJe5H3r+UuTfW4ZgbI3l2uGMgSz6Yu
NukcZdgtU0nUpfxrT7b1ZVsBwsQYDYHdJgTF+VX9mwij+1fhlS+e0uK9nk4/5Moi
MdOGX81xypZvyPSKVHS0gvXRPj3gpwdU22R++oQrEBVJbyF45XtDWu1aRGAXzvQ7
057yA1cOiqp0UB+YmHYQTxZIboW19KW+mX32+7Fsa6t4Pz+16OHUtdunc0wiMA5X
Nx3QMhqGPf/88sM0m3/eni07HidfD6eQf3W+O1GOuATE4JFxs9DZvBVfvTFEB/pk
2T7wmPgTLXlha7R3AEzpneX4mCpHahJFxSatFdinbuzM29wYJxFTpRAoc6Tx+PDo
4DyqKkFMIDAoIbV7kKKpm3Zc2joMOXr3vMtb27f0zZwDqwl4lCaVuBAfhy3wpCtA
Nq4NwLNqecH8D7EkEbTaxzkNLRhSfssneoBENbsPD+f7R2WQ0Thiwu+OMwzjxisn
sefbCnqqtZaieUtbPj6a/DGj1SYmbRKHquiBvdKIuvq6lqOEb/PRPjbCPjKE4gve
oSRaECtoKLR+6cje5Gaam/b3cauco9SJjlrasw69FFv2lHek2dDWqaevL4Ialt/K
Q3RBiOhfOXIIBNcMh+9YgtVVdgxOyAk83cPGv8a53kPedylYUgymT62Gp7uvtPg6
4ne2Uf3K5byP5a871w3Ac9wOi2/Tur3XMQ+usCOpnatzXqtqZe6W+EW4MnMPEpAp
0KEPVo9FRZUk8vH2+KIfSwncJa8eKgwYL2sPh1n+g9/OB3gmaednzqMMTrolIgxA
0xjxL61CpkYCGrx49c1sqf3slpGK9XkEq8GDO21c0E66jsWsdlFMK5YzTrEn17/k
XZQVb4G9HNtM2UPJKcbav4/cdltJo/zNOTDxqvNm9efX4bkobdYpZHz6tN7hre4/
ovmTIsH0+sMBIhibcEWolsGQy2BVdenHkE4xyJxz6Ru0CnGiXLKxFipIW6zxDZ21
aatVzfzGfVwth8g72K9G5NXSZLDWTLrzrNXM6ZPseB9CNKKbIZ4DbNSauydY1CnY
3J/phQ2vvmUJBDe/yCo+NvxiG3oW86Ld/viBmuU0eCmpdQRN1IP37O2rlKqrtk3w
bdyjwunseXYJXAIMLm69jTA0EPm0qkZAepQEZk4DXHr2cAu2FYyJwJYUU5Feaguk
VIlVsNfNte+TtY0jjQgCMKcM+PABmvn4tL6J9KwSDI+yRB4vEKLZ28hx5iJk7P1a
QuSEYVX+27dEyHdMqBL5iiXM6OS86Xv/iSunhx7q14HBv+XiahukbWOgxTmMtnIf
SjMiQH8FSR1/XnkbxmihP8XlEB0+Fmbb/vZ9gU4AFRXpn4IkTpaJQUTdDq3A2fuz
o6/qN/tJZUUfSDFIoa95opbAeNJCGKdrGHvwiriv1aH7isLueMN+0xfp9CSrhvVb
cYZaE2FC/x7GMubyQjjvylBPWZk7jz5RGYb+5ar0ZpVOkNtg1/rANlsEEY2xyeS2
2itHalftfYv7xEFzHTlCoSf96ydcanbEEF+/lhaFzVOuG0ZfsM8XnkJ2IiYV69/t
OfLS+gIAL/xfPstb9CgjgNsc2Ors2HkaVAmo78xoAmfLCrl9oVPylb1+Bg6i0kVV
sBeR2qTVyJ1pmw5ErJ34IQ2Pws3t+qBehfdxQBwZFU0kyg4ly63NqLo5049PuX7Y
AnB0PT4k7vt1vCSkphmWdDQr4KdyWotht4iuV0PPMd137WtJdl871TI/AhDhgPYy
63GOEuzmeh0LBgiSXgftw9tjeQIFpEGIz1LTyzUkB8auqj7HMMawn0V2tcIBr+/a
XM9bunUzs7VSzljyYKZvIRp1hrAzp5STaGriKCut7BW4zZrbisfL6o4iIYaZRNFi
2HG2hUo1C+n79dEwwSMR2wSp6hSYxm8LfSkZ12SLKlU0kN52V9T+z2cEL6NqD8Fc
FQUL3/Az53a/ngN9eHdIqnV7xxRq56UfAHYwO2osIYrrbO5nk49n3nL+Y2PraAo6
R/fKjdu2+wDQS27Ne+cGR15IR2CK6nZwOqcmwaDyup7PAbdYfHVGQAINKuG1bCyP
YXwC5dVyCrCIHWQjBkdqC9zdgbNL+6e7pYQXPunFh/gBgGMpd5PFKiOnj++4smkN
QBqh6bAM5xyg+tKtFFoVp97CatosdNBmTheKvrKBA5voneSE20rSLdAncMeeACEp
PPd/M3S0MoWqvOYLNKDhOV4j/edgQIoSrw3FNsiVdfUA1BCZ73fU6Ol1FvcWG4H3
YKiIRudacauyjR7ebn3PDNj8l56mZNaWAl5UM1//v6ayMoGf+WiCfDjnBmqXqGjb
Fqk2nUL9bZd0dgX/Dfhfja5mTsF8tGKIXVC7pz1pqRONunJ2Dv7BrRWoV50q7u9J
KIud/VjlQRukrz8r92BV4l8zoACxrxHil1ieBXSQ0HNnYOuf3xzOAhjyRC9y0Sot
G8pAeJyT8A+B68F/7q6y+di8l0TI0Ob/mNQuDAQoRNvZU3hvfRilQBeOjajI7vYr
27a0CV2viXMzRBynVKjyfrZ1HrDBYMrEG6ZeQTm5JC3GsGG5kgayYyqc3KlWV2eX
1THw7Cd9yQi7aoyg22wZzpMeX9sEjxhF7UKJmjFp61rYzHm2VOcJCzOf0JJK4Ahw
9iidvvw0IKVQI9qqcIf5NTMCHa9dtoJB4CQs98Gx3xtWcrkFpGrLtTX+Y5M+9Af3
c9QRud3Gf9SjmYXlFK05MJTmj//Nq6Y8BPQhDzF3CgVgc0mbCRIYWf5GH4ltZ64w
OLzfHYAmxddqu3Xoc+s9Yd1bpYrnTvrIRsSlzXr40KxRuq6aCopXef/ZOBg8Sv1T
b/9fQtCDeGiJFFS/YL1rHnOEph4dBzTdLCRTEcA0zf9aQFZXuIb9xTd19LtJCKqd
gm3t90/Ch2IqY2aNd4GxtLSK11HIl7Iww9gs9ARDmTTCl7hR5rdFvfddXsXExVfk
BhCy2yDHaJfYRk9WqcFJd8CbtC1/ZJEP3Bi9NBNfXAzkxGdo7m0jW7PvgsS1v8fm
hIZNIodXI0i6ZaNt0U73cdcLfwsUz97Qhy7TxapF/QZPeDzC9omZXPr/KCNPglHe
uSdowC3XFpLNWBOXKnH1Sx3ipJFPquMyaT3r5L/gYI8KoJ7yFrPmwVoThoGszs4S
BBtXrTDFZj6Bm6R1IfaXzzC70M16nlDwDvhRfutNdpG78Kkq69ZL6p105doU8yhS
+5XM9LA0OrGhq4BARrp//rtnteD/f79BVKLXFT1l9vRCkPw8r+YmLjOyJdsRsx+3
LMG6mMIoacRgl8zc1dgQ5p/3/Q60rOwBUGBfE1W9NOe/GNMU4I3qO8sc6I9WHdU2
EepCxkD9iwRxBY9MGnnPMtlKl4v7PIETBJY4Qk4vVyAI0WYpn2dBVly20qAE0G2A
PIgDrnhwn/pnFwjGOxUBvdsy9ncwgmkAipM4oevEa2aH8THkLXwpFKn+1UoxIdVL
DJ1QM4C+wlST8IWPSSeVDo/mCZ/ZXCsHQ0MiB0tazaPA6jSk8C3GMk5971oCWMOb
S51fWz+t2KcnAEi1WwiBRrKuflgq75qKUzLu0HBC+HuDjBqe57oCPgghD9Ekq1nr
l177Q2WMfCOsaZ1T23a2unFlihv9cheG82QQblPcalGL4lkS5W+TGu1TfPt06scG
sc8N5DpR5lMC9tAyDCvYgP26tsm33TN9JE8HOZbXXNzjnVUpBXZFGTGCE1iG8I1z
Jm7kqGQHtR/nqnIe4Yyb4zp0MJMvuelSohjc/5+45BMS5ubjkcyyulq+JGbZq4KH
s0iUmhNtGHU4Iumz/OILlLgZYaS4P/dlwLyMPip5k8OGEBi0XNUVPcs5Tl61DxwN
uZa8BBXaZy5ArLdWAaTxp9xGOAiQpAMsh6w3rfYcOFGGwaXH1ixpjhcOGVssjx1X
8iw8156U9dKarI+9a8tfWbjmmJA5NsYqugPljo87pfJ1Io7yMrW41CPS9dqcwiw8
/42EZRoEjsmcDoHXCCIR4BJEaOY2rXl87ZxVgjzqM8LCgQ778QL+MRAfjs52rj3E
wInOS8guOfTTyCHt7y4cPGElFkq0wQEd0vFjdHRuf4pCrXURVwsAu1xMYqFfE3jn
SuXG3CFirycOA2Qih4guQ2Dx7E+32sjGlzn1InQlBXyjw0ysoOeFoR0+CcdM6sW4
5mGjHeJYezzd6tsEDNMjmfldy07MjxbWQ208bMQ4sVsTPYgbdM/i5lPmiFD0yW3Q
F+wIXGfxkRW/VYFFx7pfk02z0/ElovR/oJ3zyEsWBVo3Efl6yCFroGN/WbvZLt03
GOeAPSNhMw7RzgOsw/rCSbq+no2Og8jqX9ql972zo8PIZ9O6PxJMqchSLki9gGI+
GKXzph6n5szvNLVessMEZiTK0ns0+cLIvYpEkZo1PKR+uApeHceyrqnBrR5OTV05
KbhtH6JrO486BvazmaeSkttCUBDMMhVjszP75ONjoagssrx2dgZX2uEZY3HPP7Yu
9mvFidWHCwzjC/8BGQiQHbX3NHcBxMqJTi/uN0tRopRHGkvP5T2gdrlTmuLSPNH6
ziMEZbAdUuWfojM9NCayGeElB9isy+IQamX3M+O8ctNrIwQU2fYev4NfIO5APeHh
fVgggtvVeJsigoQf2dmcIk0Y34cX0EconQeyXatC0HtBfTz34LkIO6uthLAus4OA
XdaFvD+qzRMHgISsXruorQuaZ3id3x7Nk3KRJqPMMrDchf6G8PupMrOH6Fc/35Bu
WEbnEQsaTwlMaTnf5M/+7fSQWGb2+xoyQWiF+6/y5mq46JMRpcANs9q34Mz/BuwP
/RQbIjEaX/E7rD0yYIGIl2rOSHTwg6K5BRLUC//+s74Qda9miPm5XcUb0MtlKbYv
kv3gJFu59BW+i6jLcN0CL/yw0a+4ELyIV5UZ5lEbnFOY6zRcBylBnQVigXASmqkc
N0xVLKQU4OywqmSw0JYdWtwMEdZpqaxO9CIO9X4CjxDmZ4E5TdoT3TBxcs5DJEUp
3Ne6lz3znfogD3PDlJireHycXvQRy5Oq3cKEC4GLuSdYdu7wUL81EzK686wD6gR8
UCoTvHO9Ugz1pg91cfg4edVcXGApuxYIOLH6H9jlHYXdgoNpnbPcjXAnfBDJgMG9
CpzPpccNG0VDqPUuaIxiiMIKR1GM/KqjoNJP7m2pUzAwojaXoDcjxC+8c8cYIaUS
pxIBDDkY4arCIfeEeURLnNt6uSIOXtwDURgQbo0NP/TgWwg0salwRS9VKP8fr76K
w6Oc11CvRldEW0TO3EKRysbchaQdoITqYfr+UXZCq7IU8O7VtV3J28LxqMdnGoFk
TEZsueaYQVSf68JOZV5aMUwEWAgiq0EPVG47EzXC/w9AariRg7b7Bgr+EEHWtq9n
Iq2MJJv/av/PG1gDcvMZSBRker1xKEwdey1P0JK9knS8ba7AqdrEHhQrwYY8Yxy1
FuEsiWmAOpmf4raJNTljxoBGquYVATlGLqHHjp1dC+xn8OQIKpGxKUohOM8fY1JN
cgo+zGmTuozlKJBgaDql0DFkMPjsZ+KjCRL/z+xEtZkRtez88hw4TSrc6snDUzLJ
/vypJ3N49yi7K27QgHwtHzxpdZ9wuD4X7UvOpyTBg4xJ2UCO6IYpHSS1VNffLiVc
LMlPCjQC2wAR3UpQRHb29iUfwdiGnR9Mx8ZyRyXAbEC1Fgsha6F+Ikvqjnasjwyw
XsJq3HjZSvOtDpVaruWpcOHf8zR8eThB6T1iMCjcDG8ovbibpB3dVe0fsoR0I5D9
tRAi+C28T6rUpMvem2EtQ3H7++VNmAXdpBKdJar5bKLv6RrYQ3jjAiaSM1k6oiEh
MLX86krLlWaEzCSu6D8duQn7BSvn2My7yXdj/+KfuQp9J6nOReeOr13SqHvSXeKg
G9vyt0SUNxcv4EA82eHEV8U5P/QW5rZfbJkawvV1unrl8I3dqWuu8hZNoNmF5zOt
xcT+fCjub55mzncIDbIiZyUuMe/pFtq2ejbY4aiy/zKnKbPUe9DWspwM1G31LXU3
MSp6wRSocuE1SUo4AmqdDXSkNuaQxpXyf+elpDFB+o0HbP0ToWVkP387zn3EQtn3
eEgGIaNRHTr4dct1iZ0e5u8nExtZv4oy3iVP9NsXL/fqrkkmP8tC59ZO951jrMmZ
82VbHU9Ax1kG2o/RRMAp2yzqeMXBxp/CNJUoXf/RmFRuso7ePBHGGZT5j6fnxuBQ
vkfKamFP8S3fUW3YJx6H8hp/FIg26YlR1GvjG9o2BTh/lZ/gip6R1jb6o+KpelWc
zGsaTfj4C8sK/AHi4Zk6auBrHfm7vmHZ8uGpRRbWOBeP1hXx6JHdcsJDGj93W0TG
0J7EWHHPENJsG1XFt7sgfoHqrJP/v1unFiTcOuJ6yEtt6qDBBrEd/zXKE1lve9hy
www5lGzuVJGI5Rlne0hbGIIY78dieRnutufqSoiiWZyWM0Cr5Le+wxi7EAd9f453
SR0yObtO2puR7nIvvg0mOCDNIS9c5xoQn5Vwm7XueHdpZmVE+wU6/VLBFELwJph5
IvzTgbVNrjGDW8ddtEfPZ8ESzS+/kz4AuDZABsuFjcwikGX6G8G90rxYBtF5Wd0U
3mUMq0B5/H51nHji+QHkOch3qu9J8wIRGDXTy+GcfjjCLx9WrhaiXzhg7q+/P3zq
zQqUN/yHoiRc+ET4Vf1CDNOdplz5AVDPRLevvy5gxCkr/zVs6ebl4n4Gt5hresG+
myIE9VjuAkiX5aALC1HPeEzuJCZVaXzmlkX80wXte3zpEaYSRWjZETB1Pcd3rcsI
tLiHw5TX4kiET8Au44Qrkz2AZjqAQOzO2hbVt+Ho0Z/uaUV8W1pOyBWnurajL3zH
7L38YnK5tVOvytv7HwUfcvad1VDK2Gv8AVx+QY+BVFcmN47bz5xztreDT0re8fSp
lNqTtPbSxUkYsji5SzthXkW9MS9RGiVBnku45F5TaYWl5RbXeTxr2V6dnpRl9uEt
vZHHlO47hY3W4gJR+Jv4cDVmRl3+4JxFgoD7q3phqFNYtNgo5MpD+Df1d9GfWw5l
5wFliZFNoQaNgf+rzU6vl6sMctHxjhTnMB8HCDtgkrouBWwyH+Vc9rYnGPdsjO4b
xkSJABymOsPXD52UrlF7EW6rRrxRW2BznMAvAgEArUUWBUj/Uqf0ABCG22LHKV63
N8iR2j6zEXQQ1Och4dqJkd8pTLQ4aRL6UYF1DVYefugaxeeiP1JxPMGmKd0AcGsU
99u+OqudlpyfoeQa3Ooxu7jAhT2SkJ/thn1XRfMy/1YJB4DcY0+m7e6QVDhDfoen
OG3jFFpGrAX8tYHLi2NZiGjyDSTVi7NA5RdI8ZTSVbUhjn9EnMj7KRLb+OF1GN69
bB8dDpi5+2gdfsZzgAZnd2cM/LlXsF3FQPDasDqqfzgbAGgAoT4t5qnVr9/OXdPA
z7sfOalOoCG/9g0Yg4cGK0JhlcQIDYbMqYm4BlW0JlZ4ToGxCToIT7UhaAaiV/U3
xmQmmoE+W0L27nDp7wTnJJs61gJuZQkBvf96XSLidknXJ5pa3oNH8sljDNdo/B1g
AeeOYbhoVhRHhUAdWK9r13Teb04OcpARq0YvyywBUWgIeI1bhApeYEx1yfDQ78Ij
9VvGqNqPlyYJHjQbTHjR9D9Xig02cPLbqzySNFRM68RhE+mgFJhf4cqscBSNmo+r
Euy2VC+d3G9O+GfSaDkEJNNVIPiEJNxmWNhCo8wWtYsaD9Pwy4I/wD76kS20nRBP
MVeFqYc41gbB7xNlC0Y43QpFa82bRLHnd1sj6AxWTknSfq79732DOs7F4J/9jHT+
p+7k0gTwahcmbSNLTmL7d5X9gvSXB9uwmKGE5an+Ey0CLE6Z9J53kAMIh0CukM9X
BS9dTElTQN+rt6732F86aiZo/fNeq3kDOMLGJY0J1hTIgGXWlJbju27Uktg3kFkJ
b2A+EDQ9KhYF8Y9HN2Uag8/0HhYBMvIaBBVwokuX4EmFjJPrdGHTGAXPwJ4sN3Nr
VFswPKpU/YCQG1wV+p3QykCIZE0JEquIkLb2ghiYI/X25glAHa8y2iTV5FogwuZg
RmC78/V2e/9iWHb8b6ouDf/bc9nmHXtfOxZiLO4RstnOKKcRUkJwDhKrZFSmwAmJ
QM16tXaB9Cg8pz1FkmMMOyZ2CIxVXkfVw6D2Ha8Pn61U7RCUVPc5BvJXdOiOgwCo
LiIN47i6TZaBAF1vjKvKaHxhRC7MgjAazODBVAefQMddE3J1Sea4FlJB/gi6WBVA
bEZ8fYOY9/4oHvEYOLtMpfnaMwcSRQ3zjWYUjoSAkrw3UyGwgFvo5eiZIEt/awfH
P5KEzb4NQtX/lj8AbJLIjZ736pPCujTTOxpp8OSBs0wx5IcP4z4NEn36adieNNeN
/FmwNaM+574t1RZ7cWNTkxb4MQRS2Vk2wmHqXwR0gEX+Pak5QKpeYLAtlO+6DGYE
5ZLo8SbUTh79MqnxJoDs2ubUa3A4rRv51bCJ8cXoFeMHLjL4Tj9QKKbIo85zFijA
lbzPYqmNqG4ghPqm6Pm9SovKWk5N7FWpkZIPc1CqvUopIi3CFr7XQvYY5IIj+k5W
D0mjhqlsTLURhFpPH7H5KO4P1qVA1eKpMrw3mmtfXm8PMpat0H7gqNUsUF2c53JY
Qlhrp8Ps49NJLEH4q6S4+i1sFG41edO4l9tFgxNj3maXTpCHQpzl/0ompSqMeIGG
jWpgPgYTdVqcu2iHl4OS/J/ZZq7CQdN+l8dCqKKcLl7xSXkWTVP96HAt8YVak+bg
CtKKS5rGXybeOT+Sb+LqwOz+6COdxDIyhmHSBZOfQPTpy6oiULIOUHd8v4ZEaNBu
j1nfWYBjAVIAwXq9mjivpfqcTokJZ/risjxdpgd0X8cx0UgjMew1BcThtmUeryr/
mU/9eBI2qXSoX+YTCsfFunJIox1tEgMeo79zRVwvvKhqO6PbjW9VwLQ6AijKLTvY
I0KwpoKPVU4O6QptLSyaFCeP9uIeDdSGFxl1UfGNotmMPqQZ6709vFVOypu6bQG0
/hj4BPGcUpJHFwZPrm44j1pxfPl4nk7W3ACsR8qyVJw9N2RMM7S3zZF8eSmox2tg
erV6FGh7hnSHJM023IR9Jpo6D0vLob8p+T0EI+uzYFG5tqx1z6ltvYpHRjse/7iq
phO5d0JRwJ/IjLQ6MBP4zNO4cyLWHM9Vpx66f035dVSrEoUXAq3Mj73HM0+8ZK7m
lWr/S+P7wHyR5DnRpbm2Hhgcc9kQMvyN3YP9N9KS3EsY8twzvEUp5aH2Uiw8mgJm
OqT+EX1O4DszHSWnl3BTbmPdpljhVR667H7mkuqPUJ4Ra7DT6Go8F5ZkIRaLpyuq
dZ+gEMwVYPzcHjL2d27+n7gIksHKL0gMhORzjPuT86N41BqGJOklXfuPbly3Sn4m
kAzJi/xq7I56DToqYrQeBPImThYii0THxxo0pV55jos0qc80/+1xp+jWY4WUeVlC
T30GEgFXOD6jGSdORhPCAHjalo0sTTmbRf5DBP23b9EjTFVpkGJYeh0chxYh0GvJ
skFXG8kUXccayzxFFPnSNABP83p3UAzF8RYSrKER278H07ESYEhiwTqiPQ6Cerk7
GBXEAr1rJGsIv9cb0Rv2KSJYAWqfRbql4RyuwdHMpzSM6u9Bq05tkjQM9i0nyaCc
BWZ03SY4tSnSAhsW7/Eo6kbUoqEWXZUsuuSkRyUrTAIG5FfAk7xCYOqO7a3usg3g
imBjublKyvccJ0dRR4vAHk6QAHSo8l3ey0uN1e4lLtT2gx8rOnNM5mkG1zhdZgTo
Mcx9RPi30mnMli9nGIjFHkAgvJVM8d0zSQDF9PKiRxQ6GCcvHNM9k5N9pPgnLdpO
uslovkgitrC62kb7/uCYU39Bmc7vZ0v+QB9QOllUJtF+ojJCDHmUQdM3QflPDzMB
tBiYZqKJxaKK8p4zHpneHTJD7mUekQjeexLlPrNXNEfVgpGhRTr7NpO37+IxszlB
cK1TdQpADlNHi+cSWMx08w0l2gtmdX9QiWaIbPIu1HfEXmBVMpv0Oc6orDWeT5eO
AydGIT69ESEmoZhMxJZmCa6OGO8681psSxMUa8qkktizVsONMmUYzkNJuT1GO4yT
iK85xiMMq1kcqROvB/UYp26n4NAkpzIrZ4UstbwxANmJWkCZKdC7bygyefG7BF5t
2OUmVKLa1wsZB04cC59LTNcbLB2ye6hxfdxoG5FRowae5by7W0dY1URfEqnTaMWy
8qO11hpNm24Ov5U69BDhDdZEWiFzQ1FIkRpSboTtpCXotL2lwBqPWImOEtz9jkzm
ietimbB/0/v52EMMcGYUFpTzV/64VtgH/3HbBPkkEkxJT45y4fuJRag9NH82n00u
4wIAgUo4hxQUGNqtVXQEFYsRrexY/WPSRWMrinUxQh1kwfwXqPmNbExbtz3UzolA
S+rBFmH2BpNZKHhNj8JNkKWj2fe3k5rTk+g6pFMT+hXIlfioe3Ik8u0/aJzDm9/2
TCSj7G0Z7I4Het7YTv34Iay0UqfvN2LqwmLaLiyhTnIgO+4pv7BqybAMvn0/12F9
oBLBCCHYUUD8i/a1QHbrDY2N4xYUWvJVSI8m70LHfbFCZw9HdO4EYnansCat05Km
bw+ygDxKHfX5y7OZOzQYuRpsB1cGspRRoKLmBeKI0gRBNT+o9zb08u41IPi5O9e7
lZfXpcat6fHHmJvkv7sbmMR8OnPq9RUAFT6x4MsvxRb48PN1wXw0Qw1ALaIdjRsX
0IcHBvpE5KWFWWG5yNTogNYPkOMTKu413Jeblge1WQRhXxB/CxddbjKfaiIANPl5
81Qdz/b0ie33mJaTP90waCjVeg+pEOcKK0NtyTus8VA9iGpQg2JuYjJKCV4t4DCW
REGkbDO9Jo3zeK+3f4iUxaiFuuMqm6PLrkBmW135kbDMaDnSJaNL20Sr4HH+Yi7v
UVj0q9sWlwlz679L6oDGJExvbRVWUfRLClwQ9GKpVD2VRXTg89hQ0rj3g8U+K6u0
IFZ5IlxgJJI+d5g3f15dFBF91L2GxBS3SN4ilh3xGqh9P/MZnSdyS369WxWNMzmb
/5uelcn5zbgm1uD78jRqFVk3Fisb/bgbsw6IaN2shkL4JVPWsNsEJKqXYk0/6v2+
SS9RnCu6hQUjP4ldANohY550BH1aJaSAN9pYxwhQ9hgsLobgYQ4O1MG2cCBmWowe
044u0o+UGocU1/MsqpHsKQhUuQIqpmkFkypTr0kFdGf6bnTyjOu8E5cNOLzzslzK
B36ubn9YAhw0i6MYvjxfJ1+I7Xx7IaOxWsFxU7eLnD1eS+SQGvT6aCFrKJZYjGHr
MaMWBAA/Cifo4QeK7NdSMZkXwfNm1wCFQZGYltgoE6VdVk5GF4NNCCUHRID+WdFn
FwT/u17E920VEV28MfF7yI/h7Ip+YmUzwWwXedoOPVSBVvwAenagLxOsG49MMDj7
jcIZAmMksJoWVIQRWqvqUxySqYrreIymAiqjbFtb55QWyFJKElKsRSKYPHuyWQo/
zhJOeaJ6+teS+MedOvSj7ZSiJPqMVHHAgOn89BPMGY3Z2nHAqLgvmimQeNCMet6P
vTuYRS8rB5MzQk+Xz5nkxeOE6XZMGA9+wBB6nx3jn/yLAzdqc2bnqyJz/miVkdyX
1wNS/5i8y7Of7+znwFxmRcCVFwu32J0qK09jTTp/K0ck/1OijVRJiquaB3Fp72fU
PjhFn737QSIwWDG6jrWu1l1+s0dTpUIpg39yfhfnkq68V7z1cELsNfN8Ysb0m3T/
dzM0wynouLhNPreg+gL1Aq58c+I3OQVaCIbV3HQ1f69d5kMdqxeH/vU/DBxVmqXd
H3K4fR8Afh6nGaF2W2tgdUKSEYrzQroBEz9o3eKmnYjeGfQkKmb6B5A3JtcPAhvq
aq00H9v2QrYMVmhwPtUGmCSvht95zuKPZKJE4KQAmFbTPfyKwh/kP7O+mrDK7rg+
mQhyKB1sgkAut/KzdltR4P/UTqP8ZRJUTt5VL/T9vS9g/sCU2RDWH0qiwnScd9QS
U/nxjCSrQehXYrnzMt6prJJebd7E5Q0N9fQ3bGY4SYHeKgJyRhId1b7wzN2KnZ/Q
biRamqCOrt9PK/CYejnNz8qbCUOBFW+7QCqgJjV4CKAvGYKc4QGt5xx028BLQgIE
n3RCNRmG1hP4cU6Kn1H8RyhRY6axmjbiPOsfHTDTEPVNeda6XuxuQZoyl/WJuChM
gDDbs5Pqkn3yKjnjl0sRd75ZbKcsQlQo3DruwTkDfOesNIbmEsnePoZ+fivP9Pq6
aWC3HYTbBRU2lDvfuMV6OxFjJOtBBlMOTY8hz9PzeuM48zDn2GauWgldsjRe/cDO
o8v32ah9lallIQ6BDx4k7VSfLpzghUNy2ukbhvzUICS3SyB9o0MXK6tVM+uNe0yK
r/uMLSgjNRUIbpCFfjHkwCzNfFj6MdrJB3f7FbgkbVornG8bCkphx/n4GHXNO15c
8Xd/ce3Cl/TuAwssBrI4BLYnc5XMB/Tudgocynv2qib6mvEw+cjvyrSHaarVVLcS
a0k8jdIX2HAwWII7McChwV6Sdg91k9S+9bHxg1H/JXVEp8Qugyx/TI2pNb8Yqs2L
qxkdeGemRWzJ/RgjTUIQwEj2MfYij/Y8lZHALdzs0boBIWTeqk2/h0vJdZfbEJTn
8YQZswXscCvEOApXAmHppjnY8AKIh4YShH7um7x/VgdG8z+1NbsbkoV5mFEfvfID
gYYR420JUckEh6VdjAIV6lQYydG4VhXihotXXRz1OfX8U0Zi1n9jW7ILO3bqkLHg
8syxBiVP14is8FaxQ0apXKyRTxyMP2nkuu/gu0KBwEU3yL15OCSBRLSQr951EfPN
aZ91eBQXylvjjDZvUS6jPE1l+arByY9OF1TBkbBdsa0tY++1shtYKWP6ltUJ1DWX
2XVvHA/3wcAyVJYytlxfaN9Gjr+mtY8zd5ESWecJHbQVwWC8G+cRjo5OR1BvJDnb
xdScp+ZG49YwEffKS+KJB1DSmeJHJRFeRZdVZrGasXKvaXlUNFatYi04mrnAfyj8
0217xxOiq0cwk6nHj9Hn+wPRF/Bk2QMViMivLJyoIhciayYK3N6P9b20L8TJeazP
JlFRYPr9wLA74YX3OlWQ3b7F0gpo2frnk++l8CSq1dLlb/uJP9J+rV9ffnY9dptd
MCtGV/Mwcj06XdgkMbo96nr+Tpz9LTyw9yxphlLntB5huATcZLSv+epRYuFKD3Xo
kXAWCz0PAol7jkHhdN+rTIXdhMDY6dJijxJVrGa8SCKlolj/785FKF58dktMq94z
hCguuWLAlGUdcjjcsi8C944xrM5QrbP9N6E/TN6scDYE8QgrAkZP8Wnc/wLykjUU
AOGGIsQ2Ooa18UxsxYr9JD+YWTNsm4n4qAYfUVNs11vl7lA3yatd7wOUfwvRU/uN
govvN/dQYSxCSi/XDfx9gDil2f7JvmLnqjfP2oG5Sd8BLrYZaItt42mMXjbc7RTY
UhRYT/2hgD98ptPfBJSM7/2OGiH3/hnVf8t80cd3ADggdH62jIdxXgVVnlPL3ZDX
lX4TAQKdLAbA3IlLjaunEMRNX7tLSyMrv1IcxzO68g5q4SpE7hpVRyTyy0aunO4A
LzilCa06dvfP2r0hSUlEadvh1UP4m+JuNxbN9+dudO3ZfaesOpuaESX6JFFMjuzK
rmDYyiw2dTEUXqLwsDMaxtXnrd/0EGF9yzriPHiAy+41Vwq9Ao8plJgp4wi800fY
hVOimmvetk9ZFuvIq/0VUbVIx6L5S2A9/AVgbu4/fJsorV5glwzXqtE0UbOzylIQ
uFG+bA3XvIWCk43isyV0RnLzTGmE3pFHdYNvvs3Kh6TSOxjH0jJ7nBnAossxsHvw
jc0u3zU094TEy2o43sPJObti/04sEQKPOw8mUCrcfF9vx4MMMCwPTejS4EBeqyke
M2jZEycr2n7F5nRA2cBprOqPycz6zoJC8lJq4yZ8lSgqfyQMOGKjk+DlVkpVd6+q
iwc/ZTNXO/e/2ZqPynTSGAffX883uZsVkIDC7WRfKhgVkEDLMVFj+gmpWcVeItVX
zTkk1qsWoKAhyBPLppDp0mURkFH4ujMeiDveSK2wuu/BY6zyc8wjQkiA27y6UUgH
h59LAsMbn1wqQZ3sbIjBs1B+2doRV2NVnTclT3OuBrNYVBizdEQ0I74Z3qQQ0fuA
tj4m/6JzuEMMf35RXjJL6vMmuWjWcvRoS7D/uHXIML0XNKdfVIhv0WmD4FchZkX9
0+HHOzWituE+lyFeaIB+wzpNEO4BiuWwGYP4boRVX2SHWnW4Z5Usz9M7l995phUo
G00vCD6JYtn1UwgoDvVKWKt8WHkZy5+gnUG+F5WKT4M9m4PP0OcrWWi+RzQcXCix
pRGJZPCURBQiXtLUuCvVinEWHvPjIHY7WHMAs03iNPOUqEoVOTn8aij8v8Pswtd3
WmLYVquvwNwD2RxGxHBTycgaybsrupeEq1JkcD5dPxDkks/WT6dnP7yLqvSA4XpV
KEosq5Sgxlnxa+EA/l/3M76y6kGkY7c9SjFuWFIcvCHIFgYdkicVlc/F+qzNVE/t
xTlquV881JrzK0rvg3G6PtuMG2cDEmmzPFnh8FcY5kW90A8fTO/l84Lo8JrI2c48
KdYsujGGfx7qTv6VP+Zws6bvslGcsWLFqG7+9SXV348MMsK6B3SVfHC/UHEy1bXn
Eq+5nxXcUeIJH+G2BnRwxZ+wqxKXHcygP6F/+sHe6sjHBvgsGq2NRX/1KDuQXkqY
8yRmzm2wItsA3T/UOL0VCbjHfZwkGWM4aDoeiqxWTPZ5NXAhS3vQqsM5ECq/smQr
iazN2VYhsBtlarxD+X3w3OYkdu5GY6eYm18DGxiIAQmG7YLJaFtACmAcr+LxIS44
Jqel6rYQt33nAfTirUV9Y56aWc4UlTUuQ48tDcDyEdks3PvysORfu/FyTKncNhNK
JQPcmuSAdXKzhaZqyuIwNqVNaJL8AQxxWvuwuDtUqeUANqFwlx+ktcOkdhN9wFvl
gj6k23c3pWM5+Amx2/+dgxxByCqR8AsC5IH3IalX6uJwqysSAXGh7+PSw8EDV9HA
VM9GplMJHdT1to6OREd+uPJKZzSSqNd9KBeR8TPe8cYORFYvzgpmy3+ZYz32DMqg
wJ75tlAVk0nsoZd7Ds1WNs52U4VBD4Wiceam4xf6y80U0cwC2ZWH3p5/Pcz27X01
nk8ERwRKGRVTpBATEJWuMZmXeitkv2HYc6UBFM4AP7UBrNCJRN+8lar0XYW5su1a
fiWL4yJmBmwQc9sFPPU1sFBb5XJDtAfZdncsG2WO028pqMKmCiFkgG1vMKf/pDZI
4PyXlGBHPSD9RcX9vnPutLPnMo7ERmPf/93m6vtAX3N5tPkxPEkLDyyWRhAycEHV
mtwbdVP2i9kFF6Q5TOKTb/H2EXSuRaaVkNORDh3q7mNu0jecQKceJv747uQ4iRoo
2R7zUj6RzZ3DoOw1Ip2QizzhcDHsC9+qf8cTrvsw4IttPyUKDZZjojsvTx+NtgMR
aj9oBOIS8dnKPEcE1mqbbjyP9nqeky+0sJrGjCRrhgr2wx8OzcxdAQNiNnXWd8rB
9Fi5qIXfoFvChx39MzoFOzLXcK8zedeLqLiwM4bR+L9+XoceUxFsTSsbO0JFmiWA
UGzPTSD/wjJ4Bm90REAo92fo3nf3sLR+FrjIEvpL2gkalWHPCCyRVAPxlwwA6Arj
og26CulKvLRE/ZuTY2FdgK8N970/wUHekhJwWK1R75IkHGvDWILt3lO/GM9u91SF
ro5QRSSyYKGkmoOIGxd+87rDpgoZs4hrjqfXgt42eUSALUuoXZEXrEGKVEIbnnA2
ZJVEVU6upYu5AoG6ypj9HTzTDMGpjsmEZiy0JyAo2O0FPYCMcnJE1RVtqlN7pBok
TfXq10daKapxwGAWV9uFBQUcZDf3dnp4Gq66f/kHnPCVLEX0ee0o4QhFuRPdNr16
QOj1YSBnnHIVGNOhUJ+1eHKItGzdwDqE0mUkxNWDSZuuPfMWrS8gaET2nU0cL1J8
egckIv1c/T1fPXNDM8UPHMm50pG6h2GS77Ga17NPkrU440M/mXun8le4Rzsg25fj
LTsJ5TdfIYQFqeLoaGvKUwlZewaKSdZu1nwBk7rwk+nBfFniHL7HfZm1G0G3wvFu
y9D/1/abiuw5tOByeuYVXz8ySIuzkAYil1mrD5HCDXvXPJ5/I1dUFLyZ8wsw/mFG
bNkSv01YdOlHFqnxWL1Sd87PFownV7gvJ7CdIrDUqsNA9gpnN189RWtx2DDQu3Ea
SdhWb2LNDtpiRAYZKoP0mEEm6IjOVkCKzJjBGGiKn/2X5k8UsbZ79qC+JEPxkIzD
9p7gx/F3lAKrfHnDvTxxotJ+gdNCykx+GzjidGMaBEuhf3we16pw4wlTmcF/RcPI
M3cXxVwZhfB1Z72IBMlmqJ1Gb838eX3BHoHbwzbPU4mi4VVVG5ReHtKh+WkovFP9
dh18yODg+N8jnAbrxxyhvKMAn7Ve+RTiVLpMdteg3/7vQo6hzKu9F7j+OXo9euq9
fp/itXcSeVph2UIq75POiysVsdGalrXhoqXRZn4aQtR5AqTtAPJknxI7nFAbP3b1
WsrwAk/pRMaZN+j4rRH3D6iaa6e6VbYUD6f3qK3m8aJRokC5qXdx41gottZEPsWL
yDASi7wZY1b7dCsqPZuINlU6JQLOHIv+7K3v8ekFFLMHxj+uywO84791OLIMKsy3
tr8NmZ4J5lHpwLUpic+Vkj6IRE0ZKhd9OonqEUJoelOo99EfgUeMEI7Tjs8c1aW8
bTbJ3PLqAgL/ZMSyKlNLgX/zQVS49V/RkUVNDSmo1cgNBSuilEv9i+0czJpWUJLi
zW4jbbdhxM+0s3Yvcg4x/SSWMhsjllAevEQ2oSSODYV7nZsZ86WjOQ34Z2Dp44w/
dk0tsCiEauoKVTXB/sW0OaBWvP+npom4ARry7lHPXPILlU0gJkvnKCjl6rSp3XRF
QxcwRgh8HHqVs0Q3asX0ZhZY6DF/49Z+v6Rt9DJ7DzYFTFTudbcpc/9D0phXAxKq
xM1Ih6mLkbBPTZi9vBXu+XPQMa98wqQCmy/XMaRcCdmMRoif0pX57YSUA+djHbpi
dA9cwjIRgjO0YxQk0/XEvS86+sUXymqSTWhsP+ekFkOfrnBdem1y4TtQG+cCFofW
x4/VoQavt5wsax0f4VWA+Oyx23ebkF0+EAg+hUUPZY1kWBxHIaIYPp3kzL9ry53F
IWwPnwoXFR+5OOrVDqMmx+us997VBKoLwv99UOSLP53MBLs0NYcisz7dC3ZbOf73
VYOM2I9RUhPq6sCGkFuJTJiOisuqWZdXiZJuFu+vq3GRHWdm4Rz5BQfIfbLf79D1
LjPDRf7l8RtkA8zii8okI5Vo5hBH/zwec0BzWfGc9KLixLg/41BPeihnJfHd+5YD
6aRTxVHHV+FvKh6tQROIFv6TveAeklC0ZsR0Yyeu9Batj0lrNdZJ3M5no+++hjop
LWZv0eeARq2JVtMSy2mA7aXT531SmiuEDHaO9bYDUJICijw9f4ZE3TSDr+qrQOSf
exz5DE36Aa7Oz9Iq0j62x+jsaH+y4cOkGuaN6UrhadOxJsw7rny0Up1jALNapGOP
kMAQ1xKDkdkhjpJa1J3UjNUgvccqMGsXvcU3z6+F975WDc5CcJwIet5niFb5kN1K
wwOFtPGuOjZEaIPlhYPKvJ4s7h7qLN+YMgW6PIVtw8DgS3JGwt0VoSx5RBO7rpC8
lLK7GCn6QhBtju23V/9khyfVfOFICR2ezxf7/MKMkjmk2XXMbFDAq4wqH0x2CwQs
D2pCCAJphlzOt+9cDpQ2aJcJHdPUq3f2Bj1C3EIlgTPbd30lXOuFmdPzouv0sPiu
Sikqx5NqVE9SN8akzhcEPFd56DBc5ZDm+mI4mq12TtFJskqU8Uc7KcOIEZY4EGtI
hDdFaZ9+hIRicGkF3JU4+DyC8oaIa9H/eeyQ042+fuYilnjQ8NUGZh/mvKSXu+Ow
HI9slwsEqqJBI3X9TVmGYhJOpRgmThNa2EhH9qNvvXbg88gvPs4Mw32oKIIyLYYQ
p8AXBMjnXyCvT19UU/n88F4SvJ28pUBixMxM+GTGJQtm6mOysxK3HoGZvmXP/Y3S
sihrW4EnDDaHiU+fiA+3akLXqUjAPoUNvI9y967RGBF4aM31Lmaq1PEr6+XHms7e
a1RBGBRT311RAW0QKrdeGk7xVQYlExxNqp4GjBo6as/73bNirae+UXjs0qb01C8I
ryJb+Yub0Q3/qDZjBK3/tKpwT1aPzum8A7x9VPXwt3UKLP0cKat7cyPAfHsx5Gbw
NXsU09R4Uf5UwMHRPkTWqMfTd1/rP/le4ZqtnX+9D3MxVsfl1nyV4VoCFYYZ388z
M0xVJQUAtCBQmBMxz6oudyOL6oUzhmuUe1Z1Jp+ZQGj32baqHhaRbVKE0G7Imt2f
/VPGPA2pN+rF1AwrKXwOkdq1mawUy3at+WlLGgtYYtloEPwet2ALcpx0qI7Nbw1D
/McdbA6h8FJznqtm2spq4b7ull2l12DGRatGT4CDalGRLigkQwr0Lt0LGsFx/acU
65oz4U0M7zJQ86jGrxKlMc6aPV0FudDIRGw7AYhgW3YPEqsolrkrnAvqOBc3FWsO
BSX4b+OtZZmhRU3ciO7EpNf+O/yRfZRxhejTOmNixsSj3QIAiyMa3PFJ3yrmjBAH
uYePbxcqqJ5tCFNMo6H7OGBfrrOz6XOl7ifT6BT5+BUghAdjXJTCveB0XEbRJf/w
7M85rjrlZHaT34de0XYYC/CmLgVe/cy3amv8i3vDmew344cAswe6lNSpVG3ZOLUx
XQpGnyZlPsi76DuBOEIqbtOU3JEmz6SsIXLLnHpZbCm/bAR3cbGEjfUEKQqMwtuV
mol11GNFopU0AiiuL51ReGKB6Wvxs0TnUlh7sWFkNnvq2kQKy2ixka+Vq8If0UER
M/hgcVrX8T6rojC8AD7DvZBeTpUgEQespkUoHlA+SSRpYI9yof4an45l8TKsXl25
AldXlLJlfrVzWrR+/Ezr44ToT2YGuB72qXRsUsXcfC5QRIzpnvAgpSxT2vzEtPmc
AQBb+g6dpvd4Ahfw8q48wzN2t+yk90lQ9KRfD3IhmRFzZm2OzafJ2D5k21pa2aDl
6ENTDcfMkqHlSBkMHRpYjHAPx/sKL422YdRCbITCfOuXzsltlbApANa0P1Uplzno
yYCfzcPRnKL9OI8xB9lNd2UKy+0gwHxXnzhtweVwQwtYLlzxeaDtuhpYWsRZ853v
zONjsyHScX9IK0aUs04VeKIwRWnRITZpfW4dM4qZs+f2TZog7F8/09Sf+1KypUEW
3+75PNgW2fwsiSlzxPuof2MJSrhwoy119hbSVTybYB7nk8SpZn/wrquDsJ+bL9iM
sbZVDdF0N5To7af/0hfu6y5xwx9LEWd1tW+zqpUHb2rMu2A2Z9J/w9S9H4eI0tPk
HSmjsk08sj+QUEqEgfaPjC8fwG+6/nClTQr+3Mc59b1oVqx5XCiHbJ9LbaPoELov
QHQuO3ba4NXYuXgDk0/jTm4/MalPPR5iEqdlnnUHxMPf7TUcOy0tEpA7tTiDjMj1
iOaTjga3N2gEfKRl2W3JelE+ICjLa9qlIPtlCutOT+Zu7Q5cRj0+qJ6i3nxALJDt
fI5ojlga8zPlBTxFO24Cmit7F+yOUydxaIdaJ0rEcOoIh9R73eFEA0erF7y/MXqP
CkOErq3ZyvRFGNbmnGLXA1G2FarkNT8hbAsJ/nlJt7s0LX9SMicZaOYM+TSN+xH+
J3ywyv3bhJvy/ct4//jszKVrg1FnCMI12lpn4Tt5xs4XtrLGuoU8gAqbQv4oi3Ap
UefQfwC0KtQGS6WZsc3ki25ar9feQrn96P7YDvxAyX4yedJW9GbnqgehseyNxlO6
ujuRzDOwcxBY9be9T1MWENkrH3kDa2Dh5nOgD8o4WEqEluwZdxc4eFAf9zhoEGhK
ZdbMTuOnTk7idOUByO5YmUNOp+NE7qv7zuH+go7okiriEb5r3f+Gdgp7gp+Mxg3J
Au7HFO5wnaczgq91gN1vggKevGEG7pYswvAV5S+GxLNR5ag5YsLpclad9yeYLED3
VBgIs/Mvt2JbINkv7Hjcja+2lw7gzI3zlnFO63qoJJ5MdBJTv0jRgnszPmm5XHEk
H6cQ8yGN0+NMousAPJGD/gJMoEVQ1DtqqzG0gdiAAw3Gfsq8mA1sFZExBq5LmNKH
WhuYYe2XVsd0JAzi4pXAqcAb9BAaMvHks/DZa1G7NoE4cAZsGEjNDukSpzS0CiNx
YXFjFosqP27tjCu03hWOfT3BJkz3edU3iAUaXsNMeAqS3dBUJnz8mxiCnJKmzn6/
CpXo3ivLfprEJqU+RLB2HuKhutqMiPvxRb9Z7Ux+stQdpx5YidGS+TgRXLV9cxRu
WnlayBtdUyxbxyEKh79ayo3MJsDplvikNHXGw2PkD9DNpiQkhKxluESodGpgO45Z
jzek7v3otkXKSG4lpuvGiYn8Fe8xlzyu5vkqt6UB1Ftw2khc9MR/HhwJyPd8UMTj
c6P7dExqlP/Q8MG8Vzhfe4qGnk9RX6c04Ran5DF/7YYdJ41qujYCp6MtBAYL2xS/
pwnLkN9AUt2S1YPdhJ+PMsVMocLqxZNIUMGU4gxZh9JQ6utpQYXErYnFKIemM6+J
zeghjphB98foAIqhjHweebyv8WBSnHiKWXqtD9Es+DUyx6wdmt/06CWX4AAmkwpz
7n/mVtmK8t59DpZMxb6HUaIFQKmaK3NOOLZxyq9hN/CbP6YvipZbAuYPkZ+paoSW
v8Nlf86xZWqGQ7meufmJQhptpnzY+DjC1C3bFmkv9nSO7DMur7HwXiGpftYg//jM
Qxsmri5y8+9QG3Zx5Egnh7Dzg/iGaAd6UJrZBEXUFec3AzLNsogwTWBjCBjuj9G0
6tHxxrYQ0I14iCsNMjagkrjinCG0g5903XUifJ0bWYhj/l63QuuajNzKwJwTBZjn
9od7y8AvPheCy9SWkv3tT0vFP+ZqrvuHhHgc1Aandc7BIf6njckFqoQ3GM96HiCE
Zl/RjD9CsElS+wCrpSx3fbzaF7jEjSYsgIQHbzF+xhdYFNG8/s6sgau7EGxiQj9L
3zCdVM3XsQ7WSd8ABsCBJ8WdnyrO+cK+Ik+zadkq64tjL6d8JOjR4TgFe+uB+GtM
4t4Og2aCF1/NQF2ioEZGWFgjkW1m/MP0NxSITtPYqXTB64F2DaolGWYZvZbaZCjz
aTb+kyH93O/gqKwVCTlFaMEthLikOuEULmimZ9+jNLEm1gtpQrW9NuyheHywke5l
UW9XTUjj3I/HXs6Cmzu+mU76TAF8NLTQBeor8OHgay4dcZaB3wfeMXfH8LQ1jMJq
EnjEvXemiiyqiC6MFPoZIdR5TcePpW5aRKXiSImqlCD4dSqvSOxiA3jrNEyt5UZB
OgfkFcBwIC1aRHhNXUe5vJG7RpATipyk1BjKjL9MXKQIY+p1wX/b4wT3G1CR+Rc8
J+UGPmOBkOQk1XptxYT5f1l0RmhAo9pQv0V1PkheAZ8b8S5nweh1qQaNGnpAFrY0
E9oxw9bhVY+C1iAvd2pLV8GAcwZICL8jevG/cIfjwomIToUJgu+iMn3TpJb/1oNY
ghTELEfBoqn3xVFy6ZPfhMO7bVQXw7/BBMbpbAUi/KywN6IpDiu6gDXgvFMXlUa7
J8Z2vGQ2a7Hl8cAW0DYzDbThn1oKgr0wo/pNN2w1p/p25XbB+AHI1NCBXAPEShrl
gqeGn4vAkA0fluu+TSe4sS1wvih8G+0p6qTQ1SJKisZ4jReWvlpMD1PWQITaKVgJ
rBjkoQaGk4lQXXmO8/eiwx02d2p3zzoGBWJULeG30/oJSX/N9W8SvBP8fne2Xyck
L5qQvj0Jkex6RvD2cMJt9GkDS4TCyHT3+oQgSLMVQLXFmzTFvyoMuPdzs+x4lvuA
ubso6AOSG4FilFwFw1fsi4qgafrQ6quGpQxyndXyEpv0djdUqQStYdZCcx3pXMZF
tzfdAxDst805uyFHvAatyWptl+DjQZhRouv/1+Kv5SItcJ3XHCUh2I1oUh928UuA
Q61M8B5uR+KUGlFc2yTXM0W+HRtf2ZHRolEiQXyQ1Rq95CZJUR3LVGAGI75tjunG
LZcF+MpFrdSRdl9iuo7I2XcipsHA3RPbXEY/7iDP3rvG5gz6VXf3iD1c3sk6mfpZ
s2HaZMpUz2Y5dIrNTlRKsNk3nbBlJMaJYD4mE1MSTNgSUDrQEfXi0YQiJiOAhVx0
Cn6qYdT8IiXSGmXix+vhcNa2OAQ1OhrDtLuEAUxJmQC4QnBaVEEFxQXfI5MpY83+
it5BAxRoVkTNu3sGSC9VwUs1MS/926hIMxRI1NgKiVqPZvd1cB1X8cmpzMX35RMX
NHJ2m+n3rhhbZ6gpQBx4Qik/OjlwU/AglNmI3uwso9azpcSaBecwdy9Avsa5gXZa
5a8WYgE+YdXESSPtmOmUL49hjf7er/tQR2Mj5Wb1wQsa1t92FdIM56JuRp8r5UfS
EstgyZ9lcvDmVdkc4Zu4LPPUKomvh7ljVTrmIzb3yws9u8Ec5h3SkuuFCQTIbLIT
n+PTqGCEQQ0uvfmeWdwJtCYYD/zzpItki3QnrIac/O2C44a8rh0Cgxvdu1C5sujN
baLNwnob12TOmYmaxzfQq+uaMx3TXmfHdlvTAhA/7RhjSY8pyS5k6nVvKV1j9i9d
LaXKmFzN5NqA6wgTMf/Lla3AQ87Jae0y3oWNrxxxeXZpACv9pSfRxoSNeX6fuFgR
mJJZje3KrGsJ3XlEJfyDwiTvrYXDy2RoaDRyESJKqraSA3wpRNYd28yeYUMdDTB+
UFHY2NYb3JbEXaIE5AWAl0SeWiKbRd0eQg4RPr1XI/owYIkeiRaNYQ7bCoGibcGD
vEAjgopmU/Rhy1Cl93XHDI8NfLdhMz4rXmNg46iPuI89EB+92xK2XYRuwBp95Doa
KwVLxmVMItAQCmTUWMPOymTPfmdRmgN/lSNCnWK4jdMqh32miFEOwWx3IY261QBQ
G/VnrPS5OxaUagvFZF/csr6zMPXoGNlYZhbAy+OB7tt3CQJEiswarF/LQVp8VCzY
k8PYyF6QpfdcQqjZFV+b6AEiU4x0jvbquQ4dLFy2Vxyo1Z02g8capp3uc3U/C/fy
q3rrWmlBxWAmaOITo8UP1lD0oirb0CevuLozyDRuzKSeaUeGi7ITYj6VdTv+l+hg
pbyoAsFvh1/kvzMM7FAqiO3UzYivADdywQgrkOXhoQUkg5866VMYvBTwZUirYIxZ
maRsvJ302loMZswtTZTSb8/UUGexC0nujVyuTxBqGyJmJZbohDL3ljICUlYjLZeW
biCQRrkzSrtM41P/N5LbGdDZrqWi/+MTE930LEjWbSxj/op9WHYu28gQLf0Bq+zr
NVLDgJHMhheXQYT7bjBh+8Zf1suAG9VybHpP99bXS8qGlqYowLE/D4GrAr+RKyKy
sVoniXfF9juSetqziBKbX5HtBSh4VuPuqwcZFwj8Nh1efvILnLdfnUDkuJzEV+qs
RdhJ8vYcRjmnhxkql0TgOep8qV1fCrQ1C8sjHJL8i6Wxq1allvLEThMKuioBqyjw
0og/Bs8BcQiClGgbfqSY8JDlqm/VSIL2SfjNCjlTFNesd9N/ip4qWkljNc6VpJqt
W0VhNZ5wkfV+na76XkqLZtfOrzYTo/0pW6yLNEhH1hFRyzMNY6C2ZuKzWdDZSstN
gOqoXImwwLK8FZ1S7t3NqIltIgyB5sXSxwIMrY4mLnpk1TuBL0SqlhiWFCof/vCj
esbfWnK1/wNhtLkP3AW3xRDa0fvEWxIh5JMvWjPPR/OJeeLV0X8gCEfwr7rQndz1
zpxglZAjKOOaYSnrGNkSmq2TZNucd9TyPRnDid+V67UkR5kj9Lr9tRQzlFYVvRsW
ng+jCOMy35VQhr80AkhbMtOnPSQ+JLeDnNr/beV7wkF8lD9V5GDylNRPJ5XNHmik
VJlsk2Ztg1Qy96a6Z9yc0dYky34yGIC2QtqfClKi+vjHqg+fdNky+a2WCSiVYGdr
vXzuQzTrlP8RsfWtE3O88eq9rZ2yr9CAQBAVqDqNzns/ims/wLdEuvmdko/cAU/a
PmklQUeIKKC7D36o1VMSLlcuJig9cECiw1Ye3AMDX49dXTKsXwaEWBpuTxOeUlyU
tqavXrY6ltYHXuiSO1gckvKbzaHArfy7LD5BY7jVXuBZYXBTos2I8HUHvxHEwW+a
1AN8hBmWCgyFzIhfSbaHg13BDUpueC7uW4os3FKT9WJMwxXv1d11NJsw+19P4+G1
wePeujMyYh8I4RhIyCKFFTs4oYKGV/vWoUDY5zhvEBiN818LZBxbpEgvt48P8wDe
vly4fWHZoa5MIoLp9qq1eiD+y0hhkRNrcj/7SEL1vDqR4mwVGJx8qAwzArIRXbsp
vb65APFmXQ9zwjfnZ6prKFAHtAxJdYnRyNToGaeGvnwHgvTJxtPONcqiFf+oKQ+D
w7xnUjdN7jmnw04fjXaRfpx58eevLeSecx8VXVU7W2jGSB1FPM9iU1NPaQw9KNOU
lioBsMQJ9mQ+xNy4LT+tSJijPQHzt4zlMjZPGOJnhDwCHfxA9c/OjPT7KmG/rxML
uhdEOU0aqUozN+iKWpZqPCLH2fiQkhmWIydnoxFndQhnI/G04lYY4aeS9CszfDCC
NxkK7hY7AZtWbysKxJ9Pmf8raPo14K3iKHh61EH7XshZw/qrNUHJDMx+mDFluKwe
yaPUh5G4feM68ATVisrBTbtJA3FM1hlkSGDImMLb5IvcbfTdZyVA6XHchjPzxEx/
ZjHegvcIZEBL/wqHrVVbKEnD2yZ4Dmk2/9okYfDZK/i90JJVESoayiUJ3vf+KShn
UtGYucvmOhgBaRq4XfYC4CAsB76IqQIqrUJVZ109xVppLa7lYvYubb7bEHAMoc1P
0nPHtPXSwVHNAhtJJ8Pd92EmOehi7SxF0PpZUnCWwlI2UrgzKqvdHyhvRwodiUGQ
1k5V8yoE6XVelLfpoJtU8rKwnN5bSRB4EUdb9I6XSIwhVL29RudHmARo0kzUm69s
AxRth7T6vs1cJHz5TCQufoHR0B6C85Psot+CiFBEIsfQJbmlXHjnXHG3pGLmM7Yz
5t0wUGjsbauby887BbLtZIgWyjeqOVBWx2sAcxod/15lIhqDJb6LLx8dCIFSQChp
/p3A86F9WuaCD5bGyP4VbuPxRZcmq5IJv7dBakRmxf0u7I+TAnwKYWzHMstut2qc
6ju3Xv+h4/gONq9OY9WXIPJ9SK7KQpR+P6aBqbkbCzrx1hKnhcK5diG8fA2rUnaf
BS8MC+AlC40s1Ke4zj9mnV62Jel49YOngqLq5XFfV+XxBnkUXXjXteT24+v8JjPc
xWQbltstUrSGMurCk5WDzhgU2dBExcOSUg3RMPMb8MKzD+4YYALJ9p8q/DsztGDO
nPqhTA+cOwTLJ8amzvEpIF0XpPJhQ0WgoWLpBrpU7vZUsG2WqStV8V5SsB5ipqcj
Nr9DPRdLScIJH1gq5fsiuW/8NC4gwoj6Bsz2z+j8CeVJcp2FTlizaccZZJ5FGwNX
xl6MG7rgZNBjJ+CSpUvtaByi5q57E4SBp5iS33aOIsFrdHH2uenM3Rrkhi6ne2JK
0NBp3ZqoxRmDHcPMWLUFNv5ZYNBHhUVhrXnrejsW7Qs5/Pei+27Gfd7bSc8QREnC
/7uiBkhe9Co35HY9/JrbuzokeMYQFZxeBETYHE0+/VgPxsKh6ZTNjS1LqFe1dDk1
yT0RXqbcKQtUf/uW1i8hqxScNGp0YZGpzRw9WDzdU3MsTDI9BK4+9/0ZmIG4PwEw
BSl++/qqYMkM551mSSxLIpH//FAMeke4FRUdbLDya80/EBl1X1wq2WbRBmFf9hhd
6tzWLqcHFeb0bOxweWtN1ODFbTLQIKCqF2ELT1jKubaDFEow5aoPdm+ktHdrsD1o
bogewXUGxAaLcJIg1KmmugPHj5OjFncDdy9fL1TVeycC0B2/2aMPHyz/z6mj1ZKb
7C9A5iqKHRMaXBlzEvYMzJOTz0oojSl0sDEdJ6SYdRQYTHN8j1LWbhyykVpYhUYS
QgizAgbK9VATaMvTSldKf6WP7t59rTas35nXATISaKazwpXtW7/d5h482Wrv8e+R
SzDwvBnmbFEfJ1hmUQYbYlXaWKXqG2ziE877MVtXetqZJOkZfaswmbBd+CaUGRiW
0c2aXPOE4QU5+S2A25vFE2N1c/fl5q/H9sy4XTNVg+PubnS7FVNkERXu1ZhuGpJd
dbdQXo7jFTGBWyJAnVvzHHPWl2n7Mlsz5tCaqMpPOxbrI4HhZqqW0NFHKa3p2aeD
/54fHxEccNfx/g+6y8LfuAiACkkFgtP7QtHJvRgAS27bjxlZ//bibfFLhuf3l+Iw
9+ILnKr/TAVMUzAQzlvfw8Ehtkrs7TP/JI0iHVLwZ759EIl/V81vYnGUeypx9/QS
IweGPdm8CJ3mMGIw40USi5uN/OOSJpHWTZuguZcERLJAtn4EP+1gJE37pEOPxU8b
36RDrwh2XOnDmmJRP5LvWS0k9d8zEP2TyWj5+SokodctQRN7a/iZSzBpqKGotCUO
PCIjnVgKtcXO/siAehRjRF2fFhkXMopdwfQSJMeKcOwy6l/7whJgUvnXWR5M5BUw
QtGCw4S+2r/9s5sKLrlWFxcpgzkjASQDbNaDb4tmu/nF4Af/WL45djKs8GtQCHMa
nBu36igchJWHJyVeKUxBcVfiLN4GkMLdRw+3WaIbwbAYsN64gR2+C9dnt5CWEnaf
3YM34LLV1kGXfVeBwFzGh+k0veEE+30FLcQ+FLPM76HXscs0emUVmtLuxKJxfCLy
vgIuV/3Q2w6E2EgO5o9bwBENS86Wg+lbuhwAU3GLIMz4V97+h+UHQHE8Nvuu3QTe
vNjlk2x9X+VW6l3Nt586XegRn8YjuU3aKmoo9gRWlMc+sqYbf/l9GHHKiUtxq4MH
29FFq0iQp8ggefENxr6T/aV99XQa7FmyNPkajmQcK+6dHhPJb20/GX0n1qQFGLvU
pv34vWbupp5ugTzEX3H6xGD3GxRGGWHecxPdGDDb6h8CsFmTvNBBhcRXz56w1neS
a/sLUfOsWtt7xPjNzKPbW/1bA3s98XPnx5zOhYjmyQyVhskudSL6uNK+2FiI6paU
WAmQr9MIoaoUrThUuKHnrwUSFCTqS9QByb7xhtg0pUj0CxH8j2L2u7nsWVxug6jb
qMjEPPa0ym/QUlvGVyoRyOSouNTRzzQdIka0ScmYoHMvtApCoIqsLdZBL79SnyWI
T4djGWvmrCWYb0+WkQdQ2zqa7ZOsxczMsi5UnSKZ46Lkaq6hW5qEzWiarG2VHRtM
GR5akbxyTCJXLVjVguHZDc/+q23TRkPsYDP8u2ZQ7nNGJZMZOb8BeIps0K9ncRKk
VtfeD15NWhYykCdQ97bOXDkj0PAygtcDqrwNfU3HmmNKuI/fQ9qRTFsgVUkRtBq9
D8fA8OJkKNSrMsk9ascLUn9r1OhCYr0z5evbGdLMnchmAjzChfQqhJhkUUT5LZdT
AIcyT2R4A6pySMuUYNQVRfgkcF5p1vMBmx9ZbZxBKrs9YimN04sp52+HNZ6XR0O+
ZHFGk6fWvtmscaruEuRvf/T/cxMETxr1/Y/EH2tWxh3qXdY0hGoOhB8RAsOg3fMm
Q/OW4GS4cjhgzZlpwudhpWIwhdcXCO92qjf4Ov/3xjh+F7TrsRt5kbupeIXLJD3m
rWekZrw8YQfrmub+5zzfBOb/BK5oGnS1jEXGBpmpfnLgepkphDDjk/leg7BLuO1I
GevR1roH2NzSmoWO8zRKK1fP3zJoV5BFouGylafFxZWG6s5nzxNevJ6U5XjZ9xqm
+8zRxyYscluaIwMzrUkTa9SVaCryfzh/lpESmLPyLI3snIS4rSNCT9Lg2slSJ2YG
RX1rgDfaUlfuTDgjryOUwNBHSvNetr5JjXcZDZhUxJrnI0sOwYXCZAh4rBrTOQxZ
SYEgzFheCVyUmHDoay40SdEYHjL4QHFqMbmX5QSPZGE1ITYHm29I9wnWutqbGJVB
O6DRMxoWRrbW0kIZwwdUhIE2YeVLCrp937k/WbVouCPL8rvqTWhqnTfyPiRb733c
Uc5IJrRAVp7GIA9H0KPHH2/zZJDBbc2FtEAkPRrwTt2KyveDRD2JWIv7vp3U9LAL
owp0KfbOAce4LMeNZy+LZvEXUJZgZ5dxoXULQ+QUj1Ix26eHqU54IKfYSPEMfof2
lDRWxuKIqx4Ss93cxhOIWsV7U6ictPQpg9sXlUgtM6yqn8TEd46afK28UZuVDM98
lKW1UgGASRuFacPAAe1tmCFDroIBLp5NV+hkGvPeMwsD5wvpeftPZMnBetWeE9t/
wa7t3HRaHkQQ5+kQY9o3fWaUQH1A/4j4W1iP51tuSI91j9x+yuepPc60YbYwbl1J
Jk5a7LIszNDz43LUcHoW4+M2G141lIa4MLkDudZIbxGrZ0OLC/uz2WI83wkjlEcU
bjGT/vrI49tEIZIyjbno/HCTWcrlhyeiMZYiqsysN9lcPr4aa0aRK2s2Rr1VoSNU
7NoW43ouIo4KTvFQkgrYdK6n3w0U1k3zCY/VMzqWI2uz4JKJOxdnQdOtl5neN1om
d0Y3s648t9qFJFa9Q8xoL+6xvX1z1d4saYzCubWZDgNRD7Yw3I0dRF51emQ+IcUj
V2gPSo0RQF9uifNXI2TFFG/pM0sX+xk+i07lRz/PbcL+Molktz8KUihCaZnyV/2z
h2uljV7jn4QE3BOdL/rbdQapEZWBrUJlXCaNurkzcl2MxSNdyNlQoVSRZkS69XZZ
G/Nj/SEnT5K4xXlYEbXNSlNLzHKiWvl6QpEkUOHs0oHuWEXc7exCD1lEPZ4Idy3J
cuWTuTBuYCG26GhQNOmvJVxUtvu303Zf/AvtiZA++Fnz/hi2rV+3DQkBbi4fEMkk
Vf8n4mx1T4WnjGtCIC8zZqICjrsVP81kpebO/6zo3vj5NmrcLYLNmXy0+m0jvRss
h7EbSzU96scpJhHtTR/ssPMfH29rV0AzV49Z6Bfsx6d/nLAJvg1V/puKDOt2l3OE
zE4Ew1mCLGhgYCaTogJoh4PQZBj+Oet5Z9a9FFQjoMPgRzJ9rbw1nppHgHPAiH8X
aWTVE++yObmJS/a2ZoWd+M5y7e4iARvhIt1gpfdIgGhU/1bLTMHeC6tkHi1HU5il
OfgcbG+JgW+2cgdoM8j5O7cMI5h512CN5b0OOA6Qf8mITdZZmuUxbef9InbcaekV
rgyKYpt8qrEDlUsTxXsdFYQOY6T6BkO3UeJIgcSoL+eoVcXEy4UOS4k+HECvLC7G
aS8//KjZs6Xrs1IkDfbowHX9XoMFdJBggGMADnSdGFfw6j7lzarqa9GTH/Yr+Oax
Jvdbs78kJKmOnkx5rFaIdE3W6tkoICQd2ULbOg4OoqEsJyrVtMCtYpCCvgMJl2Zq
O8v9Kqm3EFAuKGxLOE43wYItW1txaaeRP+tw7nl2PPzs9cBjV8ea2sJJuJYAk1cd
a93VgYXVJ2FDJGk5cQJW3JfSu0aEMbM80436sLpb346ICBCUSfBt8kAcK8Po6+KQ
eh9BTEM8nw11sR1ZGfP0ntWVszXaChSkzoEsyPIZKdtn9wCgzpZBlqvc3GpWjUr7
GNb2i/pNlKqr00vVQO+s99OemDP7h9dZJo9ygMr5mdzy02Dtau7Usu5uHl6HPbtV
QoNqhDLS+EBvWojM1jujGFAP+VJmn4YR9HzrNilu/5UWTent4nMpXVDT4got2zxh
DhZdF9VN+oZ+JhhqBGJnhuIEwzuX7H32o//rmEWGVHSD8Adz3dz7CiUvpmiUM2Ww
SNkiusFZQRPMVlaP0G58I+ul+KKr1GUdwMap9VfLyhTOcnm7zxfhZ11svrSN7hT9
0uOQ30vqwDo6OEPdoZjG5YEu7/UBriXGwcuGi4IPzjYv+ppoyBMsz9A667tGwWcT
gp6OopQoVkQcB208g7jmYSPY5T80z0/nuHakY3+PUsk4djI3asq0k/rqyuM6tSze
Z4hFBVl5lhay8bLledqpgec2bgFU/W8VYbZ+cjT7bN+24EftZnZw2YnC5x88OBsE
Gf5fg7pCjVtDqA7SUgjh3u3uEx43PT/YGcNg/WDavuSxLWtLbYxispNS/spErWA4
+/UQUT8Ae+Io7kWHbCpkQJjdiZW+IUS7IYLN0s6UZYqK3AIzP+cGuRbV4bUtk8Yy
ccDlxV0hrOQnZer4xfy6QYQz0uiPr2HEcWWEEyK+WsM5DlQvj2DlA9yP1DnM4J9K
7wz7K2RvAErlB1lnGYAMUO4nheCqfsjc91F6DbXbQkRgXyZiSYezW2RdI2wo3KXL
hQENYTSBhrGeOpUXSqYt7+gUEUA/zd2oZGJH5jdgy8DuVwM+DhJSF4RrmkIHUsxR
tc+qfXwmYVDacTbI1cvM9AFlHLJ0hI/o4Khc9hGGFnX1kPnQmVfwjZ42XWmUvaSj
GUCJEGHHa+aGVhodA0HeSrYCi5/rpN+msrvcSj1eiJGTcd9H7B2gVmDaD7HleGOS
Cy0azK2iAoTN8vmdrwGC1qyx/IDclCRcfMECpmGOONGwnT+ePdASbSBmMFXmhu+G
ft0XNaOSGrGMP9Se4ugYnaIQOjWRMwcVLVq8Uav3IRIf/CsGxOJ1cgyHkrA2H+86
3HleOptqQ62S9/dhdzYGRNHdHh5bCCyc0XFHOmhHv090nd6+A94nUBfNEuXdqjK3
icI7/xy9FXxWEvaJ7Ywf+GrTLUXwwKmC9T81jqFt7c705BeDKUH4hgVo2Lew43HZ
ghFN3nqcrrZnfXJ6CLQRG6l523MqMF7kWAnCnc4G50bfX26XWMO4hti0fC8HPYSq
FKgqX8uxbav7z54/mZUJGsHKQpsR+RXgG209A3E7Ll6uBUdwrYqR8Tpxz0Fev+aW
xhZ/EdkZP/gu5aWlBfusURPmCFuRz7XsP+30cD4bwZHQRWohdAEIbTmNVdP8AJgm
1C4kcxztoZON81kd0kwXhFZRs68qjMYdAhvm05LVNtZ3We/NGgT6UUcSDrfMszCc
+ZoW81RR1FbWhqSoz/hijt6kaRLL7FzipD4nihbRmmFDDpDm8EMZ8i5pcN7O/f3e
wwsxB0EZFe4O2pK0/LrYjNWtH2IliuZY3Hl2c7ZqnXNPsYAgKNQHTXQVY+KdBSr7
tsmpFBP1pd6Fcc0xF8WDFEANd4GxB3sWVHwH4+i3tMOfV9SQFwiH4R13ItDlOXUH
HjU27BNWatpz7h6fxQRXDFT5n6ipyqaora8Ob+Q0GUGezZyJtqA7XWD+CcDXhStW
RjokeonrpaNepwgoqvFIcRlVfL//C3wcWi/OHRIGClOOdx1zzhIffD8T94naZUyN
ySNkngLmpIXCXS0Tt7SY6Xvwj2DHsBazhn4ceAJh0btgGqSZBIx0d0Qrn4j1iBhm
+9PB+yf5CB/hcdC3M00ebiRj1/2bsVMo7Qr58R6pDV9MZHs1hfsjN7vNoaNhhy9N
AI6et8e8MYxofR14eN4uZMdfsf8prKVz43TYIGGJrVx/W2BKN1cnuoSrCf6rf/Hr
oyyrP8fuVo9wZQJ9/1e3xX66/FeQcWy6J09nQpeLwxfSIE0H2QK6xPQ0LSs5qiFR
Q3GjonUiOmFNQI7OFW8mlt7jrPgnKfIVdXX5cYuCNl+v2iJiTlhpL7wv5fky6WEE
6NBDL2cHIusguevx0Vfo/arlAcqh5xb2gvnfWzwzSWJyL3nG/5d7kN3678lI3RIS
E4p9XR7wZ+Sy6YUZ2UjSKvR6bUhPSeDElXFmngBX6fw2KithsND2v1MitJQxH4Tg
lICEPeVoz2VWf7oSU69z8BN7i+AJE/cDD/ponr00ww9bR6MEmrYAhKbZDVx0oLxZ
iA6U8dNHMYfS6sdOWUcI216HKpGyadiUGQTUOpW+gMcWkIv1MQExN4NEKN7mQ1DE
P7/HNbK4+7pRzxpFwzmbbc0v0bEeUzAQfiRaiCXDvU1T9yaFe+8dRyFPxiuzpbi7
zlBIOWW/cfvx2yceYkEwA5qW3IoJEA6cK3UvLto8Cn60+AbFbGIJHMnoEdwfxefu
j2Mb2nFQqDMSvuv8+e1oy7B3t+mxAU2LqVjjvjjpdCohYnOkaYsgYKu/UkO/UEUk
bBCk5w40xlKpmXnyAcNmHEObE4DLSXfs+Wn+qzp4bqLCoH9x40UQo370UyCMyGn0
KwpT/QllnX4j881qRpYIihLvpvLbTWIv2uvBnXJJDufswFlsv/FHXPGD86tubjdP
Il2LjKTEYVnb7QHf2yxuYiDY+/DX3CoGsBFZ+lc5tNhkD4meTxqjBLyEy4VOguqI
ZWRljySPPVEM/jwBJLiJkVvkClHfJtxPdhSS1yJfoc7jkCuFMDx0WHLu+NHyL0Ar
rgqgfu8t4pUOCeD28dwElfnE3DlH1yTFlZfFGFC5/zvcIH9JYXMt3w3/kGsEzYIF
27gcuvz35hn+ShPivcm8nMgGxT6Yt4nRSGRmJnHEzKTb6ayGYoGh8oqCd+SZZnJ5
R6kE2yMGZLA7YzvJQB+TAGuMDwLqRAVqKHC/QAvYN9T9dwOvhpEKNEP8cAlNGo9V
ShX0yYI01koBTrUts9evha6OyvKKN0H5DEOGlrZa4vn4LK4reOcIBT/Hc4pNuNKS
0q647k3Sh2qTxQY+Znw9FOgqvHrzHeqmHKIy3ILc+kvmLQT+Hq1wg8eja769u11u
osyXu2A8q0rncVChkSiqzehiTxSkqjBkj2SSjoPtaO04bKK8rrCb96VuOIp9A5ev
gO1imvJxJLEMPMtaNhtucXv2um21sjifzhcr2VpfoSAYx8LZm6IBBNKuRrB+Cv+g
ok/Z7bRr2kzW32se/D8EMyYvmL5frij4Ny5NKncW0/NMy0THuaMYBPn+6UqmEhZB
ED8e5pce1Eo49/OdTfgfY52DHNiwxBqTlEzLFaNSamwzK98mM5mpSHLCDlH/XoSq
JuN0XWyl7Ao6mQA0KOzQpiqEvS8tFbRCmjaiVp9WZMGhvOOOEKGtzUMCJhslQxup
oAYVFZI2xtHMotygw0MQOaYg/bOgSjPKmNTQK+bDo7sydo4OrgCoMP6y0ww7iTST
2t58Mh6UbJVG9YVdgVZNXvXQZE+/aovKEnLe0AyuL+MOyo/774uSyCUPjtsv1Ukt
GjvbjvhuL5A5v1SzXgQsTkOr1Ilxo/4068LRzwFJn0lUKJ0mB18gKMJ+3OlvsGbj
nkermRA/Y7I20ACUkjaSibB4Jpod0EP2ro/AOyMectRmdwebhixjyy4EFy1D8HfB
3rNYaaUyrKzO59bVxour6wWoAzvTVSQfiwLec3V4cebH8hwOU2VrqURwWwZ5r8yq
/C/V9Hy5Gj/XvU8RwJjzl0YnI4bGQGk44jTS7tons9q74xvDPeYGNoGnDdY9M4Ir
9oL3NgzchLZSCo9XRtyywG6j6P2RxToDFlzZP/QkUtX1Oni1UuX+9eCQuzvtjIjb
ilg2wQJfdprLRSELBfsQpOdHMxm3npORJYGxKDdGvke6qFbn+xPly0dFiS4eZxDw
3l4EjV4p8ukKcykm50qqJRF4XRkmjsGHrXwzrlUoHxRHuycu0n7yheBCKzAtji1A
fAVDftwgJAf04VGGnGvujzTAlpfWJ88XrhHonm186fRx+8or2mUliB1TioPsASCt
QrZhVaQWhluUYnBogC5YeJQvcn4WIvpoqIZvyBMU/U+ucMZIMFlgQCL7slSV3f+k
nAJTJ85lC5ISHo4lGy7YUvXWPb2DOw7x02I4bX2g86uz3yRr8wzxDDTgdEW5/UH3
BdmZQz0StmQQnFyXb0VLw26Boj2YmietXA+lSXXSCutjWPBWno5qoEtK/WVQ+4Gx
+md0c7z4sHEpGXNDNR2X8g+prrT7dSAKW3njGo5U/LUsf10dLwfH0UQqxWcrPboW
pFcPj01n/BfDv1uBivavGwANIvdW5KjgQs/w6cKSr9lp3cuVcVjFuwQH4VDlpAS8
6EA5WvXhgFGr6f5tJ2S+tJ1g4wPWyjUKcS9mDYydTbZGlBpZBW1r5yzuynAcxIyj
C0vFS297NOFTXSJ9D39gjOG8b5ozc5WcUW0Br7uFyXC7Gz6aJtj9gGEPivbom6oT
CMQ5Bvg7o5Lb82R3EvFqAoJi2+N3FHWR0kFFlHbeY31QQQk7XetZQNooMFUUo62r
5ZhcOI/LWqXLC4pNdvMIK1d0RST+ZstYWadCCnwy+Ei7uIn4Jr0erGoyM6zSe4BT
SVPMniDPqIf7HKzvbKdsNeEDtdIoUM4H6IynaQ/AQcViWRx4jGcjwZnvHbhN7yN6
OiZwLuaTd4iCxhUV818W4tKhcqIaNMOg4d9F7fIvWaIjgea9uJMKhwv6nND/lt7x
ShZSZcvJCXvfOXxwzShTNjtd08tyYGRGMkA1sbz4PE+w6Pg1TfqIkTPIJIqXCf6b
fccDJ7jYJYnzm90IDF4cmB2zm4KAaNnGEmW+id1j7GTtYkyQQ09xPZZf7TpRUIC/
BWEq1YZ3wtVig0cDlcyUPP7zUty5yZarX0oeI4HO3vCfdCa1KoBv80uEGvUui3wT
noXJdTuaK1wU8ulmNTCdqwF9qOSZsRvhnfVXgyQ+MpHEAsM+ZQin97jaG/J4fsBY
LAEMQ3H9mrCuodB/k28Fsj/Lf4GXtAr1zMQWiby9PnOWMNdEwU08c7Ca/q8SW+wk
rOgGoMaYtpNFtAqhvHUMJu19fzEcGTz1D1fqKXemsrs5gJjXoCeksmZ82eBj0sVk
ExVowyTwsoa4V/+V5gg02Vz6Vw2qWThX2W3MVfMZpa50pA6TK/mORO150KYdSHln
f0oQWi8i4qcwEnhPxhRpQqr2HtZz7CQ6B09TqFmpDuI2ceZWNLHxzbWMCPQ1QML5
u6iviSW56miMhUgLJQG2hI0X9E9D83uMy5GQzpHrUDomRU/3d9TpFJ0to8Cp7Ben
oSQCWDvm+vep668+EcH2xkdWDdZuaqHR2ufReVAAoCuLcyzaAVDyNAljmFDcR5jp
eQs30iU0PhAhql+KieNxEkJJ00PQiKmDKLpt95y/oOv/aWdWBHST44DKg47okuAj
nucX1BlNRx/Jm8XOjmhZQgWiKU4alof0d03ufGhYSdXH0yu71XaZyRzIwFANB2kj
GO2sk77w2Iykpab6EhGy/nL45GyUrPAcnZeM2UvSMnoaQDLegA6kYpxMe0W/61aM
a3QdfAesdr7yJqLWXO+mFC6+kUQtmZ10T4oqxb2yOCdPJvLL+7OqYrbk+XuvTbep
pqECBrEe6iTNeXOu8oNq/NaLiMl9M5oLPLkhr/A+HPy404WHLvlIHwV0QTHHT9Zz
ElOOl/LlKdUCsszwfPRtpRCg+4UAKHKhiuGE0j6tGPyOiaOXZ8InEEz1iKx7tl1O
+Nd39qiA64viN8XM4BVjS1XRYdA8xxkjm0jQx/cLDw0/IJIUMV1+SIZ9e8AoicHR
MgCTKJI9V4xuoFQNF9/AkxuaayMFmYyB44RhrEz3kT7Y/b/a82CxxvPB9nOQjjXy
Lloum5TR9p6g963Ida8haHRtAuvAOPd7G/Zo/to4ylbd+rBWDmMQb747lpsMntkw
Zj1wslZls0a0khz0S/22FMpizqDtpFjB0UotvAIdLsDbZkd+lJBPMv9rwEK7WZLc
cQBA7byhGlOGFOlvQE8ykCcGndqPOz0BNGooYIJ68CUg0zmOZVjdR98nFgudC68Z
4GYvTU9uP4jAw6VWaO14LnpcEzloLytuMGL38gkUfvCp3JyP+thKVkDVbdHOM1re
/QCPERK9taTCQGMSm1pvhJ1FxcJBhESPjxV/Fdbf353ZAPCB9TcWQCFVeKeQmhbp
x4xwRE2dItQcm2BV7ctyezYFCvZ29FSVL1QjfMY/7AWP+t5Ir0/6ng40JXg3K76a
4vGH+MSM00vAx+Bwbzp5KxwmRUQlAYL0pBp055oAsZC0qQN2Q4CPm//e5za8AhXU
rbP4XtvvRMvvCuS8TAAe8ki7SURy2YTg+n7Oo8GjsC4TL9qt9HWZ2LmBtBwk1gWP
aZ6bBZeCGZS4EdDXIPJnVfcyQG3dNIsi03lPGv+lGshR1P8blgborZ2sI0jPXHa8
mMuhgClIO/CZ45W5U2wxgBTZNVNU9LePKtGDZcUDEgb80YlwtvY0wdqY1tNqKT31
PWdL66VLMpAZxGB6gCxLthTXO5WaFV6aqub7SK7NsW1bJM/slRhRJJRfmaI+0vLX
lBXGmHLjbxba9y2Nsl6P0xhqqQVR6qN0HbigxMq+uEHV/X2Umyig2PXRReJ6MaKQ
e+aiRQ4/LLBTT6AVXb4RtSvg6+U/QnTE3TFxR84gojQzOhYjusJ2hVcSo62XVbBh
QrExzQeF7/XZJcWIEWle+kXlzQ/87CbUnMDrIwSbbTUFczpmbQCjFvUJQ1W8cAdV
zPrReRiU29INUOrMdWgF4cRPLr8CU7lJiovYWxGp+/0/ryDbOMwcgYOq/xxbnxP6
gU7yrzHB+ViZp88p9GmUAU5ZCxKD+FznjKQA60wQYmq4VE8f+FisVnPKbLu37Ys6
loTycHmBCGkh3rHSuhrPCCSzEyAO4U88z5X3Wqr+TiZ3qGnhCwvD3HEAqs8AuJam
JZGv858KdFFaMLltLh4xZEL+ltUm2gjD/zbn5BPeLyaybTJJ2ITUNCnQ88Rf94Bv
7NTuMKQtT/E0vCM7DFIOG8CEI3xJB27w59NzXpLjn1UeoEbNUlcpffS+/QCoeVjF
FyonpprJBmA8LlpqtSWIFz8OJykYmCDiD+t7tcJjRbSy3ExL3mkbiZxTdO9qWnej
an3mjB0sed279ffZXCioAkJGvN6eRlgn6Lg2+rm+8lbDq9d/zFkEfKvQ5HfS08Qi
tlnA1PvTmdaU4y2uCoGFy6dD28fa/LKGXckys9kTET0PdeSbHaoNKdaRqtDr4QWK
h7WpZJUfMu78rHp0U3THDIT/18KcA9wy+xb4vIcWOhlJRSfgtI4aZD6A6h3PKwn+
KotAK+c30wiHW/ujfAuNwWungyD1EoI1UxJb2W+TNFJMd1JE7Sgp6qbtHeEIQgCd
CmkZbL531S/UK9yWK3LVck+8c/xtNejsVUtNOyFHCXzoFLilq5xFc6lB16iFESv2
TZP70i01vInr8t61KjKe+tYemyWA3DtbYtEKmFhZgLABvIu7HQvHJnflrQzo1wuG
5bdvUcr/YHQ0nUG01vw2cWtHJyWWOd4hl3HIaws85mzTffk5oHH01HFuMBDsQgfz
68adreotceWGziBUmMJWURx80aEFoY11u2ZxOkcNwJsQFtnUPLjDQInuoVvjrGpa
jHxN/kxMJunBCxJaGkHgieyDi83LN8bDxv9xVy/BT0NJ3nbqsCvlT8KD0PwhFLFr
WlXS6d49bd0gsiHc5gz0MlPApUbsU3/SdYME5Am578o5+HqyYTk5bgAjFsGmJ5vL
TtxfSr6tMo2aNaL4Ctdt+06kDKpW9uzBUA+RuQVurvwFZSjRZ0JHWTuqh5MipydO
Dp0uKliU0g5qM67vRQXczdw50uViJzmi92XMbT6wmLOP4duj3c4kaWd1xo5YuCUK
ltcV3EC1tkbzwxgH9Lk7Pec2dYZqGZoXW5t5RsvxXqAiKSpnJ8ktSVSqTW/cNrit
F+GfYorq52uG6qTtZXNAJBb70yjFWShzCwLAl9wdX6q2RnRpzcOD2JGMYTdAkSpq
eIU4jPBruhbPfwVhGpFoesXvxDA1XszXUEvrQNm8Hc+rP2QTYu1uMfGfU1+wx4Yt
HMUjHQ/755lYUzPJhTUS3+qqTWH4UOhpL7Mi1UrWHNnfQpz69XcLJe9wsCxB6joK
6Xg3jq+sYaigqP0ISKitlHMSIRmyKTkVoyD7NKn4vxzcEqOdU+aO4Hi9H7eMbzGm
s2A6C9zpbJds139/leBqaOH90k6uHSKTirB+GgU2+O2mV4bb8hu+uqoi46s3DJ56
cYT4tM18OLVUQs9n4FPDFhqeKuWL8CXVM4CfsQFLPh6JRBwfovBnh0C+LL7m7Vo3
wOMEKcfm0sREPWlNS6naTv+K6sG3wgdtZKd1B2VUZRJGY3b0MHtDoJ+hMI9VMqBy
0lbM7OmDyzMrgELPjexZUDUQpMY/pGqKOu+krjDHgrgkJSBD1+NH+awJBuchTcjp
G+lj2ljNHjc0haZdS4+1sqQZ8BZrdOBGkfrcn1Du12QW93XnHjhVtsJq9N8VNicQ
7YlGa3t3o3Bkzhywnys0rC6w19Y5WZFj4l38ssMeTLVl62iyJ8xGcO7MHsfrmx3J
o2GAA7Fb6h2wfMR83uYzlHQS0Lycteua/idpdeA7FOypMZoWtfQEc9m/IEMCeW7G
vKc3CGxrG573iEXRx5/F9C2uEhjfhNUwjEzI5vpBgfCGNieO9AVXanerQPezrQEZ
CDM1YZAA3Z9fzblrK5piZeWOGfCXHR7f2JlYH7EtvH09FlhqQbOnRf0PVZ72YSi9
g5R1i8rGzRJla5sc6VOsIvzxVp/iwWt/uK40mzxOd7rTN2Ig95rTh2LVMOTz8sIi
+OY0MhRUtgSZwsZ+L2CoMPptAcC7tG7qMj7atqHcebLzceUr8LR/9sXHpVviB1lS
SOHmELQMgJIpRoh3SEeZeLlUtm2a3SwZRg/pvVfU/YfmpFjYIv0xsgYa3TNFNlHk
OmUwrXyNhdtb3DiqEgbDmb/PXgZ1in+n5LSqWyuggTSSIicShFIsPC7EJ5LkdIPo
CbWsHdoQCdGNaLek6ONjJ3R0y5E5XTtyj73WC3WfZFkm705F/Yu0q4xry5sF/c3y
CX4l5j9MIPlwM6yYDPzq4hGVI2sw+nXgLYthzScYou0laIspoNEYV47D+jUFzRKB
pIwQ8gw/datUzb+cJ4RR2ARlMZdvg0CcwcEIhY8SLJvhZaNxZ1FTPxGuRbvWFtkx
tK0Mwn0QGO1A16Uhdk/mjK9Efa9bXWhVhuc97VbZgNugN29mRnbAbkK56t7Q1rWm
5SYhDHNl7lCSMFrIXk1Llv5AhY17YWeYT5/IpTGZr5JndLez6Cy3xFqIlJfuRG3M
i4Sf2wLnL2kpRApJd3JrD9X0CypnpKAfD5++oAr4OLsUqL7dtWKREmLLx2Iv9YY9
Qv280K1lUd1KVGyQXSjJiaayjl/MIUG68c3Ui+fmom2S4JJmNTK5QtoNfogHx13F
YAnHZDyltbrGK7142LOa+/e0PujiNT7l1D91dRydAyVettNfxHu0O5YTVQxqT1hb
l8tfvt5FGKvthLkx8dcGd0xIbISAHA8psYbhtrZ4nRa1WNjv77jY9oY2MHVPtgU3
PjHsH7Cc9wXPcx94tRdysImk7MkDv35CtKkj918Efv5+DwU52PMa8/07U/hwNFtX
UCic81r/Rs6o7targ/iDxJDQ2kiVHHH0FwGzkUhF2uB4hx14vLVW8CIGfd+BTcMH
wDl8Vl1djO1LeLpJyjaZYAA/ZzEQnipmu4gMm1lm3S/o5TZPeM+Wmd8TEtRxJdaM
PGBia2xOXzj7oXXQZWpukFc/82BXYdz8MG/TRE+gNTQy6U1esOD7wb/4CMa3230E
Nf4K3FeUlccD5LThbpHdXAIkw3kvAu7Yl7sm+cACcaStnD338Iz/Nv4NeAgLdVmU
zCNbmGvsdMs8OGGchTeSQUWOkF9vbsgxPKL7lrKkRshCZBRvqORS6GpdS3uBAcOQ
nNY2n00EkhOUzP3U4eEuI5ZTlom5KdpDvdDrzvhorlt5hxNVBbsmD2Wm0mT3ovmt
0MfJJm2VrMQxq6ddj2VTnvDF7rjA3FI6YM1h8YRphjQjWzRoZF6/d17DL97Djg5p
cZx7EhMhZnenvW0uyNpIx1YSLswqursOT1Se3wYrS1+9cWkpW0wHegAqBwWci0cD
1lg8pQg/lRxyhehtDx0U0t6aUijjuTEjI7SdK0dVwtNrzEkFQiuN2wcndYmaGXyS
0Ar5dM8Z67AsYIRtgvIbBEumLbYhMZPtoTH5GYZRVY9x5BBv2kYeFnEhVfbqDwvM
B5s/5WL1uOE9nzlJfU297MTJpHnSfd45WJ9qRNUiV+Ltk1BK17+mAsdYqazzc9gy
E3KpK/ANTMPIT5NiwJkspDA11BLwa6H3A8J7fSyvDl/y11E1NGXkigso7IdMOFep
FKRIz9RfcthllM1jBni8UA3YdP2Zy+mYg9Eo0vyIUwW8uCMNSn0fz/DU70zWCjd6
1zVy0I5d5/jwHGdJ5RqdVrKtm1beFbAi3VHhz/3HWj850dFFMvPa4K7VHTwfQn5L
gRo2k5caX4F+eYGaAgIBy+thu1T3zGna/trW8HNfdUSjofti9k/YlU6yLuC4oaw3
GgyHqVW1Tz3sfXyXw+KMS7gN33eSIHfMMOs2WZibWzATYUGUJTH6LhuZ9R/ZBuAI
J/zyhZ2AIW81my6L+BKAwMaW5hbXpE48qX2xmjDDnw8szGtO9fRNYkLW6pIb6kI0
BqMtEmTcUA0kbDepLJH160KNaQp7k5T0Cwv+Nl+POapeX615MwivcllbW/PTSez9
Atp3UIhNWhNYVWo6XwrDk1lKu3NQclemWDbdSFlzkrRSFe2dqcFPcHBhFJkJE4ea
MDt05n9a91Z30qpoJUZNL23oRmZcpZ6jUvO2bDppJG30xGH1H3tSbfp3Z2PjIBrX
SRIhxmiAr2aItA/OF3hnLgyBdKSgEDKpA0fW8yGcl0YDfjliNJfHP7bK2j9gMnWv
runaEErz8axRcPWFBcJXgO15p4mQMr9g69GPGKI/oOgkUT/zwKA2W0tWOAeugZR+
I48hajEgRr97snjO6+BxyUJqvJN8kKP9dDse3TEZSj91VNt5XuBXmbY7zdTtGbtg
hY+D2FRyrPD44iKfN8odr2pk15bHWVHt6OumFvKHrM9H8Zh4OUTWW+UbvS9J0c6B
RKPSX3b77rbdBvaPT9LphjubeKI/qt3N2qblkKjr2VfmTwZ/52AnXoikEfchBver
WJE9SB3vWtFHzqESCv92JyQR//h/KheQOpc0gG3hKCZNl+RX/A0Au/bzokkMMTRh
XaKhhXehTtZWXtAjWGSFIvga0F7KEu1v5QJvFuTnGpN1nfsjK6IYuGUFpEL+MJa2
UL20WFodmkbVTO96fsVJtRwB8fJTcsN04hPQ8W/QVzAAqNrdat6HMf8KxnrS1Li2
D4dyR2qtZPh9JN/VwKfzoRTGqbeSThX2tm2oBuDx3nkKl9v7I6JqJ+E924uoO0A5
PG1ZoXQDPBnoi1Y+VQvWOUUgnq/pP7CD+4DPigdeZIU/KXJAg6AK7WJyRGb13851
5FxdgiJoHKO5O0Xdz4qbxin8DT8PhfnY2YP4c2tH2mypEci2iOxS5I9kzsw6SC2D
Y1+rIlKiAP1+YOUhoxTDCYUhWiIoENJO69m/B30D5V59ncuCpI79qEGaPEseX4lF
cKrv3HLgaibicV5vGxlJho8LbiBXNWh49Vjl2yMKORT6jbJigo70pr7QShCupTNS
gW7f/eML31oP9NnrwjTK9JuDqlFt6ixwdsrKm9glfKkuR5SV8ZxHm2UQEY7ZiHvk
dmJHGTdDIiKyuy+cPj3ytoG69jLXWwSZj4zeaEdxIcX/PxetBJCJ7VFlhLr6F3G8
FmpF6cAuDTQxajUmzssmaOw3RMwY/08+h0Dzg1u7uY5SiffCqnNCTQyP3fVCIfpQ
8cnw4X3Ga68Ir26nRwippeICK0Y1t3LrTJL860SP38kQAU3AKLHSYVoRE1kdDHR9
Lv3VpTtbOozRZbujEQC2xY8BDnywxetSnqD3P/wJPcvJdPZ/DBFHQdv/p4qLFsKb
qMFSezBjGfF5h8iOyfKNHWsHcE0G/vArbksSCU0npHNVzKjiTGm08bXNpIE5lz5J
RFY2hy07EZ/M3twNQT3R97CGb3vpAp5XJ+LUmoU9GUHNU5/t4Zs5ZaGRYNJ3CwQx
low7x4ZWs2uOPXsndAugKQ/FG+eEp5MMUFXEY5F64ZOzTtdLrCO4RTl6nhAEYEHd
1pI4R5LpdaSjec4qlKv8xCkUUO2dQK/2YD5o87cBkrEu+c4ci5GSBj5caSaGcTUf
2sng9vAAO3IUtEkqZuhgTqBJVHbSqy/hMP7paw+AaGsTRsQou3J04wPrxVlUF4zQ
dlhrlhCNq2IAc/UrrfHbjQidSDJ4OCIahlM8g+edXhGmH5ZVfcWwrlefBPEFdnFP
T3jU6PYwDzYEjC8ZiUG4LlkU3apuJ67bjKnzHD5bz6umxZ9aexMMzk0LM+bZ79uO
GTp/+nHMqyIMOGYkEsyBhvGX5YC1UUT7mCz5U94FEYEH2/ideFIzw0sQsiG6I9L6
hbdzBuAbUilp7zDRibKew7CrPbc0SI7UPX4acNgR8QMczKprNyDo8VwledUUaSs8
51LFfxp/AnE5/WML7HGOio1buHbdAlvAswny7n8dpsnnmz02FqFEpJGPiY8CbgWS
mwBIs9vN1Cg++zIJHYzTDS6Cfas8XecQkVswssnc3lLqlnL196i+M2tCAw6Rngoz
u2qhhz4m1rUUODTZ03SUqBE0xCpVRRPCVs1ezFNqM5/NYBL8utT2c+91qIxhUMxy
7CGRoLgelomhqq5tDZi7NWnrsZU3E3eFfTDbrBi1sSkTlL0NJ+71i+/uZJy9sBNk
TK0d1pgOH/b2uXjDoJizdW7gyZBK0X/7Ohxvmfig67p/2VVxd1yA3XfCPchiYVIW
i+LhhZRdtJa5mWoIM/62lSuVfkNa6zXzliv0g5nJawl7aRaS1bzW0MQsmOW4WroA
020nF+lIqbpBxGw0eXDyexHblBNfN8Xk+PvJTqxho45w91GYD8CDvOZl6BXvkz9s
FLE8vhShguNtDAlKARcBocM1B3z4ApqBwjs85S5Sa5bl1UB+hAJcYZpW+feZKx73
1MhhgDqZEImj+r8i4+7BONygM6mgU0jgxIUm5vgsbOUhilkVWzyELjlbyfrpNgZA
VgJWGtjBoKpHLu25OUxbB8Mv17F37ZhNnZpw6PezwT71BVdw2RnwUew1LMy4lcsT
iRupCzELxuwZTf3OpGpi6W7GrSK3FxWqfF/oX4oZ/4rKinGuStBsloAecak5G/l3
63RFzx6+VWrdQoy5kgMKmuA0YNkgpQThyAyyUlVKVKb6EgkxO5qVjvUyiFn7qt9I
YOM9xZNMQ7iCZJHl4hRr14P651AwEi38A14V8yJTh67bJ9Ei0R2noObbFfMUgSOC
zi1CDn2Bjvj48DKcVRpbCpMzafWJ30IdS+8iS3L1/ugV1z0o6vV1kBnUcjtmexi6
YfsTd48wYOzsWhm5wRWB+8L6Hr4O5XjTOPvpIJOGf94bqkIMhJDAhbB/VIYwqQIa
vCIZDK+XVkl+jVZc69Jiz0Opqwu1XbaoQKsvJFZlbV4j17TQtHwkiQsFloUATojr
IEcFuILidHahgxpTqxWcE5g5szJXHu1dIHMB4uraiTAUgk8tcajxeSPbGnOxJuK9
oY5TABeNeRr/ezVNunJs4L6q7XZ2QVa/8pQMQRFNIvoO100LKvetVgW+z+ucbGH3
/nYXWweSInNbeSMiOUNWNJkLdPvVjfU2INd932/Fptt1B7evCrfN76YQqa1iAXA5
vORFlM0Gr1rsX3l/YhyVj2Gbw0nVnv8Ajp1vkdcyFgFsN/cTBasqkF+NVL2m6VbO
AoFc1yiWrHuTaIgXDGiC+VyGM63A8nZOI/mvpwRbGiMd9EIcPMTBDs0lDzUBE8c1
Fz0VmLwKGgRn/j0QRDRyL/Va9GfCiQwWGumwWCPy7Tf+6sktBsqXtVJMUriEzM+y
NeDHgzYWUvZ5LaIl3FUIyne/udYrOG2rTuQvhEJg5TvHhhgdvGP4+wN2ptHrGny4
4jodSVpB60JbIphbwBukmYcqcALyVf92KeVo+90Nn2oP9FIF8s+TzWzHHBraUHjz
kEqKestfhTSCEbHhDPQFMyJCljgkqbgCpAuJlj5UrWH8GzSWMrh6QQXuO3+5VMN3
Cmg0oGSCv2GDwttADLtQ63rUpOnRbOido2GXgf7ZihmLchOuHJjJQxclFqWZLqXn
KVz87xJori06/6Lwqfdkvlsnzfics9FRKbWiBnPYVrRqDlQDzt3KgkpSvDfU413u
xOGnwG7Bu6/v9vVNvB0ugIkwojBptcMa3CeTvFzZ73PXMAry0LTohFdO/9rm4U+B
KmynBgi3/B6kymsAcItmS9H6XlG9GV2m+sWwHytuhjAAitiGYAgYDWVzVj5tQ+LD
GmOGmdK0tOTltYbI47nlRM+/vQQen7/bnW65e5reZrI/4YiHxQwBZXoe8QnqYivs
iwfbQZJ/LjqdAWyDEVz0ReqEsRBCqite39tzGjE62sZKUotClG1tx2x+UPwgTA7f
JqhXDLYFmgzWPARF6/9t2ftK3iqqZMJ8+v9opsRAIN3Hi4jX7WAqAJxBuqQ2WToE
UlZf3/YPghmC0GQDXAfpOWsOpZQhJk9w0s0Ts/xBGB5nnzdaSWivgx0/1roiEPdZ
x9c8wERqBwfpoB5BszYj2zBTXciA55A5Ynssne3r/d3Lu18q/CsJGpTMrtVhFuvF
TtlBNQUw/pKX/NkDPLrcN2mZ4/wCb8Nfd+gW8Kjz1REiam95hgHZ5o1Iwxxw69zE
CKIMF6tLEkAsZknZXyDjhS28uloQG5aLdJ8HBkwNdFCZK4Y70uQgBKny5aiw6YFa
CXBDnY7h5j+8sLe2GmGv6ZANAbbWuKF/+g7VEAsJ/Eex5sDJCwJZlD6GjQSTESlp
/y6+rj00blZHPnz/XQQjZHphEFNOd6S0ZW1ONuenkZq100nnA4l06D+Ok/AXSoIy
M4t6sxq3cN0MS1CtusxOaaXDENgevFvyD6Jigwdrx+esklykmtwylFk3wNDd1yKt
IJpZrxrJYVU0jyxXMlW9p2I2D0EZysFtevbiqZCJGydThKb39zvHgo4/kvWWMGbP
4Ug8lGfEaQCL7La6EKUP5vNEi2msNSlxm1GHWvqhOWK1qY3fk7ijkVSCgZXypvW7
JOL6dB59/hiwVq4XbwVhw0ExMmeMwyKR5rYdh+CU2Z6TA/vTij9kiobKx/zgD6sy
N82e214Olkfi5JMZ4irV+iDhuFC6HuqZPRg9pRvnZgWBpa6FReOvT6WFuZHrQURa
9g2siGsEFpIZQwuxfdQIYsR144/U+jwrPt8Zj30sqO0eMh8A8ITkmUEqbwUC5m+z
uJtpIzoSBi948XW9aO+l8QYlPuEnymVRjLcchk3HjqNeyXdw3M/9a3h+0TAo2H9y
1G3vADd9RgxJ4ytNYaGImp5HbKM/M3+t70EAWyR1R/Z/dnNp6hTUr8mWx0/UZCNO
TzblTLDl4+niwfWq/7qvQMOX0g2jVoL5BW+jY4mF2wZwqbFTfLjyqr0QG6KesYaK
QVpJ/98fj0nyX7mVzOYRP/Iyp6Lhi/F1h+nwgdXxf5QONy1gZ/Envado94T83BS9
hERN3SSzBocAtDf8nCb/S7iDOPHsRDvRG/5a7gqE5zgqGJkLeoOGSTh2gBR/rL6Q
L8HaonhRmcOB5z2U2kC9DhwM0ZAiuDV5hZQTR8vhJrGcJ6WzAwbVaftImVhJjSq/
PoDONliDuQ38thoINUkP4XEN2YqoPhvIuROtOGHFp5ZMA+eylOErBxlgj4zrtRcz
2TtmE9i3dg9vzLh5NKedXM3cRxkACTMPxetIooZZZVodRMlXxSpbsrooUGfee2oT
mWOJGDRwJ9TMI2nnBcAz5Y14zu/L8WYgXUL8dqVHwnmkHERET0HjWsqijE3P0qnv
Ak5OLdw2byfw/DsSlFTlbUPsd6S5X18h70nlhvnaCQLHWUjSaPBNB14bYLeC7JGm
i9Huk8oj9Y2MsCE4ubA4lvpsZ5Qt03mqLwwPhCIg65ura9MfH44RvviyYWqo3fGK
LhoaXFfQoi0fEort5IYTjnEPTr7Fdem+8uCeDKOuyN+F95fdUATma/zNwxO9Q6G5
Gi+aoJXLgIjDAHb9FsJg35ogwQSpHjdgA7G/7iv9CSh4/OgNF52ECATjodFqzxa1
K+CKtWfsQ4rU51dKD99wjbTdtzm2mixV6YzhmGnmhSiL8DR8ihsP3vP1WnpjDw8f
J4kN6B3hNvc1k6Son02a2ZGlS9qOCFusLOkNLTSDcsfdgdNQZLG/hWj3RhJU4M/o
9LFclI5UBgJGqTWFURl7HxoYqxvDP5/9HAwV47yAsSCmK5L8ANp9CFg02hDwXuCN
UaJYyA+nXxGqm7C9BVQp+y+nKs30l40ei413rRTyxl7Ix+g5nwH6Tbyd4knlwYrY
ULAwRgl2PsN3RhGnuUWpj2BOm9XpcoMe+bH3Fp7eRi9iyBXL2sW/jLP6R/fVlWKz
OsWFGT893KZNBOjchpkiWuIKq3nsGnYH7PHcI2oLtdMZ/Kbet0SRWRqqDIt8oWYq
e+e6AMGw27toist6KE0tvxkiBXdKtaoThiAFFikx5GBRksZQX1InhXrJkXKwZenj
J6N0a/GdSEX+B0W1v1R4uNUlu16xhin37Z5wDRxgUdRHTY5rjvryHf5SrFBvBW+f
P9jZOsZ47TV5Gt3Ku3xYcG+ehN5JbDdFNXLoOZnDvLDpU2bjjnPCe0vyWoH6sRMp
o4sp1iVSHWEyb5xiMiRd/hzfLXkTCxxFAeHoHF9/YKpCh5a4+EyITFsGwzBBCsZO
Bp+R+XVf9oKv0C3AW7B13gNXnVdL0haU3+lPhSF2ocVx9vOeUd4TrZYI114NraIT
gLuzSsOm77SHhB+iALnwAxXlzKe5h+NwnyULFUAcCmKzkXZeGYhim5ziqzT7wzkQ
LSH5FX9/v1WmGO7GDEoDhe2tUHO+D8Sk+anXTBzhrH+M/rY0QzQqeAEWm2dl7jAm
HeULUXLqkz6nVPlg7uAD+MbnD4l64k8cuD1BeFXja6PqekCX5OQIXgs/eAET5ErG
t6LCj3efVEIDjvNl4SBAMW3BooP7/gvtw7oO5hkGl07NjsgjGJ8QF0PnSmYPyg1y
Cv68vhxge9Ftyqs7ktSiyqkFEkmyWBKG0OxQwTv9l1AldZY6on9FoIFCfPQsJIPV
YnvItV6STlyVP7tjfOX22pQQx+L5GEZvDmAdJzAuKdU/0l3tL07zqSZ0hvqD1jNx
7ng6dS2qBW8XFimqJZdUXeZ4KlLYfm/T/mphVjeikYfqmmIoe+fAeUY2/6lzqSm7
eT+0iNIG9bCWGZisB5Rk8PXZFABxR94uQDAuQHnro2SEM9DXuYmzZPYGent1VtGs
PXbdJUNR9KkcUyFjV1tnE7ZWsydBG6xlhjoH7NmCyeurt35xD/JLzo+nMAJ22aoj
ydWBV0/a/qxQ8fSX1mddGWMVfhLI2+MfhL14K1kD7yrLi7gKYOhVAs5q7IIDazyC
cpZ1yZtuBq1dftK/uGz2kLTD8EehKI/wfVhKO1q99TVN0dGIdCR/C2kayBupHcaI
G/cQhubg/tL3Ixlk6MXq8+NNgRhoJnrEgDHQP7XhdQnpNOCa62zo12gOYHv6sMjx
f+RD2r429+NivQZ2f9XTpDHHOzRimf657YMynh4AEdcuBfYU6zoPzhsCspgiTmE+
G9/GOmpst9uDcDTu4fN7X99XBmwrKsCQLrY2j6LLdjzoGNBn7C3xXGdaFzmiwJs2
jSzmlIz6Z3Qjqip+96Q56lIYPjbqviN/fKgUoSLRj7QaoQZ1nuwdbkPGdkDUjpYo
CSZuljiGRqtookfEtJk4O9uh3699FiGUc90PtMFsRZQTSPBbBBm6hrnXa8ABVDAD
PultNzEnoxm5ukvJay7f4siGPQ4WIoI4doqdXZ6+51nTtLFWxJqBIzroJqp7qhkE
KMkObw1o8B5J8kSsSE9Yv7ZuQpG577lVD5rvx4b0H8ZmAt3SOaKjRI3rRr0T3z9k
Zg+MAhA8A+6RtC3lVqCgWn5CV4ItajzdxUjGxnlHalWhCZmPYn5DEqnrxxAoEoBq
T8I3DtCzsF89xonq839DfCMc2uju41Lp2lYbIpvLDW1TVj7gdnRyNA8eQqLJThe7
+6xXYajDh/32CUZWWWfzg8ZrDkfR3bPdjwoLmEzPYzR7r1M0rbkNQm22ynezUR7L
U83IBb/rsKTuhT1b2pVMuFx/1Lff3hRRhtPKylAdDz0fA6FQNK5B81LhYGWxnRRY
bY4CjN/sAYr8jmGEXdoEXuEDxgAmT98+NTJO9jdJwXBCrlrlm+tzZvO86GQtjV/U
XGYCLVkR1U+4jaDtnY46tIa5zkqMDIJghdJzasRaSof+wUOK5mlwO1Fp6EhZeyYu
MWwZDhwLtAk+S5u7siXtzPSpZVr15xQHDpZ2U8IN/fFAFTjwmVjd0K70VGarPfLx
D7golQL4nCkGlXNYXm5HKlsytCJV4x/0YtRf1WS31ewMw6R92DPxEO5wM+vF5JC9
zs0+5zxrLROI0nuv4Ogryiqz7OjXZ+GMQYlrDKlWcnQHrLXwN8OAePsdR+dlU6Hd
NQl1A7usSonNAHyJkQYPm0+wvpliq+8D6vmMnu/0bm/kLUboqS7p5TerF+3Tz9jl
+Wjdm4gHp8Cxhx5EMVyNvCI+8v72o1t/aMNcRbpXiyjgiAo8HMGUbgELnXvWZuVO
n8DR5+Ul9gx689zZ6BN1tHvfzH/dhotoiqo7TGbk7KWCOTZCdfvaWF7f3oZjACQj
1JMtSiuFeoZZMQ4ZJSFePd9YZMYntNn0b0LGBSQjW0AS5z1OAGyCy20N6st4yyGJ
/LYmBsqbevu5Cnu6/V4pBe79WkfX86ku/DdCCTeVupKsdpSaok/l1QQW3Q0wke8x
4BDgs9W05+4QPfkG0R/2xNwK19SwIjQM1SIJpll/2A8wy6JhJmbzmOB+cmvSJJoh
xmB8qNljFPW75MHWhRVz+PJVeBybJ9V+2qAcrYG8KjKKXQ3X4Fv4Wd6xWF+RNO4o
OIRu9jFUbMrcSzAad2HQVMDU5hwzL4pXzWRcUQm0K3MTtfWT3ptcIjJjHfT5Iuiv
etHFApqyUtBGhXqlNh/uIVj3U9Sq8fsz1BTIJEdSOnirxceXYzYoeist/wjk9uD7
x+LTLDGRZvmP2/+XA7bQ4W+Z4zW+KzbbGc6B9iXe1KRAFDyRGypp6z9KxGwPc681
41IBMWgDsom4lk3fIU5p+k3U4pLeTqsDk/xTmXYn4BC5IcJIVQgSOyx03THIyyZ4
mQ5Qexch7e9d7n9lv0OCC5km1GHjoHtNfK+A8zQRUGAUQqNtPuw7dcBIKdiPAX60
P++Mx/1HNc0pDN7IXKwQQ3+FbvkloHpvDKLOsxc1+S1vE6KjHlGlpft0riT7Buda
L5sXkSjCiWYUrDON7wilcYYetn/PeehLo8+YRY+1fVpWEmuEO7hQ6XSeXM247CeX
eI0hC6Rct/Us/OnLZ1lKceh4dAUlv0kHKcGtYTXJhxKkebCK3apidkVwcIgaCKP3
ynuFgolqLfz85/7hGkVBtj34iU/z9yQsdkhFucbyE4C6FkUmMY5SGGWV29eRUrH2
AkbrPV+obg/v8p06VTCqhShf1qLrmgy+b0Cb/pRPapBtsrDQvTxaVG64x2SZZtQk
8f3EVWLQm1Wb1UFf0jdDP6Uj+uAKQxhvSI1MRxV+fMXIk3GRLhWpcBmwJc/7oaji
vnfMrr4r/5+cM/0x+3p5CcLhusn1HvkeeCTUbFmLi/oGM1z/MQmeeM4DwiQgzGY/
xNwbMGrvpXiKqiTJg7uuiiQxS9KasPLX+/tjbzy7GQ4qPqrY9Se6iF78P3zkdh1F
G/Z4akZglr6qO8qRuxiaP0lcEDhIcgN6uueOejnkerMdr8m7xORv5Bv2N9hXJ+kc
Gr0w8Ll83+DBFuYdPu162sK3AX9LYp435sRIAjBc/H0cY+5AzmbD30FgWvebODyI
vXrWXKZ6JpdBezQuEzUBJ2eV15xsFVpFBDVVR+PA2Ao7onwaO/EU2llT0y0g61ii
CwiIWMM4kNlOu47NZKVqtgf2qGadVesOjxEujAiHhoY3Ko7uQE77agA2bEZMGlyv
xDKmFYvn4PFzDDT4YJOA6St60l1rY9TyVEIMs7zzdTQtvPrxafyTMI3nQTF2TuGC
tM8cJ1sCmNZLx/aqmqO6sHyS/QLLes9JlRkC2v6pvfUeLfYlaz2B/4kRcxGW22jm
uawAmYkGFE4AKkbT5HrUxWg2bHlF+EESyeDiRZTXW/UEpqeCm1Y/bZcstJ/pheqn
NBhX9mh5MMy662LYFX4Ylmw20FJJ90R6nN1L5ymLm5oecYqSBHf1SVmDHhGmSpnV
dKO9AOLHbgS2Nfs5P1lAI8KCpkaghphDw7RbGSsan2kSRZsKpW6/diI7WKNk1S7f
Pl6rxNi2PnPWlX92MGmLPKJ41f0qdaX1fMedFTLlmPRFMWB5pRaLF7teW2rnGzBT
DIUECqGLirVOqSiWWKAelT3TA+svhzh5wT9ClZdyOZX/5+GZgj0RasEeDmgrzpFo
BgVpYN+fZh+PAPVZD5ADnUazBH8QcxBzWkO0rn50OXM48hQJbH3cmIFUPUwYa/W7
Gn8wkO8m9D32JaQ8nIDgW4jdxdUART2yR2tU3S5ppY93TQnK5yHCQZok1WDRiXrN
i1R4T8BHW+iItZqY9hrSqc8B8oLzrzItGse3OdvwEkw7P4lUJSpZp8nQZqSTplHp
Nns4dJFXe9pLNVENgzJTcot5X0l17xcOtuFDGVAyOIMfOfDPkJ5dlA3aFMqkqf4f
bZgiNZuPaHNXLtp4A81UD9OqUVa3MtSf0ohhuDMK+HdkbdUED2VhngNa3lKSCeGH
LPagJ+OzJuTClTduJ2wg8PudAtd2PcfU9CSUmIUIaCd+G1c9/u4ZMPWqX7W4RO8J
Ew1uinyYh2crywFXRGS1SG9s+or6+wKiMlBM40lH9ryPOytx03inqog022QYBguE
SUYpOGw+nuE6G5gX/QmM9f1TKwiX/mydmZR24zPVwqzwatweXkiBSzN/Al2faNoI
5fDFhtDtitBX6wLe/PZgElcKCLxMVyCmyYEi6LScFUmabHTi29m5SzYbAxQrFneQ
erCuvo0dE/FUh80g4IARyzTR5DBVQOpbQdT0VjuJmI7hlkyBm37K0RV1L8kH3AEw
Kyw+JynlwRFGgy81h4X49tOfe0xNQsLNYUh0s+eqQ6ms85I5fAxC2vrzJQaQZN1t
qVjnBXdJFrIQNowAcNvw0Cb/Mr4vA/Ay7+SQS4iDyQtog1GYBIX+IiU5Z/pixanJ
8SGyFA0hiIsuGn3XrMY2jBzCq7IfQWYgETKS0W7D2pfNFrhWQBKfOQHS6IzVULGS
bAWJ7TlVwWN7Bbtj4KKfLYbLmTh7FfOq7Mf3ZpZouL8nGPCRyNx0wyQzuVxpOqRW
2ymnhLg6tZc7a9PIZhWKB2f6VrHfGTultPeX1OkeAEKlFr4MTNOCkCh+WZTXpSsQ
VuwvmO9bhtp/lo07+sDAd4jB9baPO9HqU7qK+fdtef76hreGRl220q0JbHznLX2B
Qph8n13KJVsu3rrN4zZin0V6ck99WeAN/RZJszHPx54Cr16QTWgBjqfWl9wqnDJN
/5D1w+kttmOFtTVdjC8c7bCsYYj7ZkzrxaPGntNBLdxTzbgmqRQ4WgBEPbVSm6aw
tTmoGp15HNwQNH4w49phDIDcPSTD28zqRrdFU0Gt4sga5vD1In/vNQCQBAw4YENy
D970ikstjtIhLhwsk4ADg8yufR9CKzb6Zu5zJsHAEn4ZakMjoE156WUmI4JDTbDY
Zy3HS1Uhiobcx4gKf30QgQQ5+//bKIPK+0T+VjPEOrXgQrhG15gkmJL6+SHmeiFh
hqchqJkuu/v9mj6hJ48SIXSe4DBuvO/w7EtzMtLKlVYcl0qKl50RoVHLTxF/4OCU
mtepUVmRr/cksJelGlO7qkSnf582gNuvhFlvY1JcuMx11okhc2Yn0ewsitQT9oVA
Pmemg0WdcfvXe5riVx0wMzjrwMJO6IJL5l+iS05He3nq6QoyhfDTuYpLH+OIi4Dq
+oh3a5FcxqTFMCbedfXaNxYs7vV4VAtRpvn7kXbOcPG/Ngdbu199EhpPStxWumRo
724Or3dvh/SiWHH7HZXoFQ5Eymxev9Qv/w3htDPABwfWKR8r7cSSC73pf9AQv/FM
UfA3Mw/F8KhviunDEIns3sY2C3Wy1ivPR92TSRXJGfZPkuMxUVo2zgFHynAW6BKO
r++Td+0bnN/YZ4QKB1EUOq3hY4OgqgdkGRobqaPIjBiHcEck+tTnnQ7mnQb56gZo
Ya7dhttTMndwtFVAH7FiDzGyDYRh1WqQiUrn4j/5CHkWiGH5wF1R6CYQMJemwkHA
VVAG4DF2We8g+ktVJOd9B3CPbRb2V8tn8hgIOQ5bdQ94aOcm7cfD9nl6yoyFlfqc
Pv4N9eZDTtGPUrwHJvK/FIQwj9mpjL/qbmEeC8lHZ7WbA00mJlPq/YYaePbHSfmm
4CRT36qr/lZXyldxNrgGVg7RM4CUCAch+REsx2F/dCJk0Kh7Ieq+3NV/LTN1fWEB
Iew/rmMJp8yWvDR8Hx28BF1EY1R+LfvLqnPICzt5K444yj7FEPbZAxhQWhdiu4e6
BNyYguXOU+va6wfZG0GYG/0ixDoTWmdeAkvGzcnrkCMR1oxuW/V6A1ur74yr9Ot+
WvUHPr+eiQehVy+w6Fi4wsBqw0qSfYiecyylXvpD3tQ/A9Jp6IEgAkmHdLr5vv3v
dG5b6P5g3dY1zxX/6gSZEYfwokF3ZaRofquqRGqYqujuJkD8dI3p6PEncAFa9Pt2
J7uAllqXXr+XvSiH3Vr5pF2pYmyOUhTTlKF9N7MhQHCAs2Q4tzrj2UjQCBz4I3eu
bOXqOaC0lmOObzoJwYFn5W/ovOmOdTHo/yWJFuu184GRWh1eGaDDEVBxQGpS0/5D
HPS04q80cWno+I41yWeaCc9ZFAQLhwWN7itMI3vrpO54T2DP9H52GA6zjfQCpshb
LZLTd02ZkNMiwi6bY2J7LHcaTiA8z03XZbpNpEEHQ8JR/oI/gZi657rtcxCNLD6s
Mg/REHSR5hLOm6Wyk8xEN55ipTXc7sLjrh6G4Msm0v3OKLwXT3vL22FTkVPJLEIA
cnSD+7GUi/drgdKMY882abSnSXis2FIQTm7E6fkwqnzqOSa1aRn2EidougCWIiCQ
6h5q3l1kWbcBKFtxfCCP1UpiyziO+BMVqEskzM45eHcM0m/Nu5ZdeQFzrDrLfaMi
Js+CxuPy1JXij+rLSdBYixjLC1RqqdkGrdgw2BtTdeyDzEz3bEYkdbBXgvwZFzRZ
IDoWExRnAXkdosR+N9jVSoBT1gAWur8IQ22tdMxIWA6CwiDE6NN7JOOKXQLGe35a
x7OS1+NJL8aTnp6E9qaSjHUtleopZ3Ixf32HCi3Eevrr2pc+yM0yL3s5orqkagw2
3DoRInIknQq9j2JDZik6C99oc4oxJvuYYDnmmn6z6ulN2Zatf5jXXxpjGIlJf+1k
hUZ/5rf4iVjeRk9D1HHSh2dk+iN8lih9jAiJZzd8eQ6iKfAWXDg/StlZyX1CzFwF
/dI/wP7T6hBCgt25XG8qOG9p8QhDKBvZlyYGjd/RcoNCRiBSaFZ8WzFrfFQhaY/X
VJEqdgMI7F/hLJSd3e4ynEdn8tSqT1iGerrXmUH8e6cQC9F2kadfSZqPGDAqz5Bc
bT9H+l5/MVbIsHuftLpYfVxAGD/dhAwsnZkEwcYeB13oq/cbi+4Urj5GCYzXFl1+
r1gmeJT+4Nh9nTCUypGGGs1uv4Olz3/mX3A8GLhqEWqEaoWEO59L4sKkvigJvfJy
WR0U72kYhtZdZFbBzZcG2N9KzMNCTUba11WBpu/q4ltA/TIQzESTrxTYfWg6Xbvr
1XUBW6n1JRyNtsBzlODlyuCqbR8/Scwq6Mu704pYw48RFS144OJdohZpCytjggm9
s2QcmLjIHODuyE/H/9mcSNlCWvzCq7t6UzXbvtT8/6bMcrmmiYAE4JEIC9FxwzXV
EkV92vUu2CW9KcNkkGaPiA+9fJVQZGVigxryayn4VcSByZfsCiBnPpJFegL3dBh3
Qj+FpJxXhxJQjbqfjbYJsKcQrosxLTL80YJJg1P/SJITAKqD87FhwbrNWXnLQoTv
L+qRuzAsN2sCuW1Sakdqpw4MVeuGNQlI/xx57McZI2wMKSuyRlC0iNti8cx7tenb
zTbOm6BCaniPhKj6eoVwHLHcToVOUVZOWerOoqIz2uiP058uULepsbJhSD+7u7U1
nzYzIDMmiCPwTpLi49TzAez8zQEMZnm6U1OwWubmJzqX8W8ljWp/2u/qAMPhP0YK
HYiTMC/r/kH/+N32O7enuBfiFVfc/ynZcM1jD5tBsDWOm+E5bNhQeVOl3ULyUNIf
41wTH4OhzGUFkjw0FT0NrZJXScqi0+H0yVd3UvBoohL8eC8aqxyRmX2Oyl8F63pY
I4ngOF4cK7gjxX8WNnSLwfa97Qt+hCRmlyQapAXR7TN/Q3y1QFVbGglziaxZBa17
Th9ZSDhMOk7uyGfte8bwNNPDh4W71Q2UDTD6ETZ/DrVlhVHoSpog8PKdB1uvt3/l
hrZRbH97ZHY4ldJBgpYeu21z7V11BHelKLvybJTtXVM06m2Y9lz89AP1b8mC4m+s
wmii448JhN0t52VQGC4Dc3FwoxipufZrsPFWyY00OmMQFm1BNxNVPz3nj6o+u4en
N+Nehi0UJduI6w0Q6/WinP36eovCqhTdhyG2XuCyXYTnvwxYyL/Ona7QFAMRiR05
O8bydrBwR1iVA3/Aowq1AB0BSfzz4qK0NmK5kk19i+mgG3Zabje4YQ2ijM+UOs3M
8bFJId8oJRV0sdggafu2x+iwcbzBRyMxAo6NFuZWxktiSwTJ+s+sZEk7HAm/jn28
P88k1CCpYAG/LXzBeKgL+TDm6qQBd8bCjdilyVfq01/S1NcTVXaRlVytNRxKswo0
1axb9HJABvyQYmp7JcErCbwYvuynEnDVeHEericRdNPAo2LQYH9b8e3zRraWYTiN
3zpQRRa+T2SuwJC/uA0GYQA191Gkav+tLT3wHP9ikta/K63est1J1v2xGlg3CT0C
vmYX8A5ibJC50gdZEuSPuYSmTj+/VdlYuYBk2+cb7KBpeXZXnMPqpLtGhWM91Y/T
Z7MtOawQKXYhipKw331QSXpew+ISvZZlg2jkTEky64fyCHGfq+vSY+woIA24XZHy
vKESUPlRW2VVFbtm3Im57N/riQJVsw8z1RxQgCeb29/gqaOXww/xQNTT//vdjLuf
mPUSGM2Oric6CK514mZBB+xQ3Uafm0sbHx+JRMh7Ny06eQqqlUSSXLSxbuipO2fB
iABjNdTtVNFTuCulhEnfnAgTq3SiKDTMs91CEkDIxqJ4QTR9Xwym2/rjTo/tMTSi
FQs3r7Y5sfOE53AtJHfDvUt7qwrN56HprpHHHA8I0bhYTmT61BpDQFib8kJmniyE
+eIlUur04EOrhXxeGSfMlIcajLJvvD3J0UUrGV8/4X9zyoCgwCvHimxRxo3ATooF
xMqt/zyMl2Qzo/b6a8yxw49KOSGta0mB8wINoJrfmNv4xakx9rShyuNpgQnfBCHR
6vA3ThTEvO6T+Q6NlVs9lO6WssAh/ukRtSscD8A106ZNGAzRBR60WY/qQ1EW8UXb
NGVW/lelwdmdBjDXXll5w0T4ldjEml2JVocIGtGkMGowHKm+ZD57xg8p9QW7b6jS
IMZn9plLwoy7x1lna2ftlElx71A4rsaNAuENiPsa7NNI9OWpJKmBGsRh+SLsXQFb
oNsxpgjraEtC0Oh8LhP77RrJ17CW/NdPzZiXPrRdnny4eer2A9E3CupIXDW84mPL
JqiL5jYWY2Fjoz45jBj23p7FVzrypW5WEuGvXUAVev4Gg3MfA6WFcWzAehmUSfaw
MEcx0+gx+/83GhYepW2ZHGOTSzc3PB1jLVow8U1FtSZNnST56Py7SXig0ltdjkiN
YCwQ1Vk/y7dpZfAV8vsbSV5DSI8liNzdu5tqFfLekwHfe9w6CLeo+fMBsxy0CIOB
38JXPi3ONROyoF+WEqxmEWcbGCY+WflOYhH6f0aCi1/kAfb4yUQYw6/tkxdMnyVd
6SISrV9A8Czu0kIk4a09NxHDiNB4yeYAzqxprZjwbLJ5ws8pw+oZccT3AifIrLqb
37jxWwKLV4dsNZ4T0kigMxWSL2OOz/l0j7keHfnb+C+tArKTtqJlCLnoiAFZJHo2
C0jsAyaCs+kxh4uzK1itj7kkCZjEvvUPzA8Q81MEaXSoenHIfn95THgK6yFZUp8R
Am9yRG47DnOVQuAcSTZk1ESLYFrZre28VoAQsA1d1K9QowzEkuupfovlM9zsu7rE
HQpT+75yAl9Mn7UVuXmlu8ht6TmaMpdu9XOkPzDHZR/GQk95tl2FMM1hQnrQ0mb+
SdYEvVk/qiGYFJChca9NSBY90ZaowW/3sGQtuM5UKQUKkxfBIETY9+mffVtCUfdV
zj42/SR07OwfDOTGFk/qYmnSsdFVwFULwrUjyqiacRynSoLvuaDQhBiRMzPOQ0k6
n82Wmkf9OUX4BfXOUrafI8jTkeiM67nLn71PTx6NFghIWoCvswBWuGvlkaIbTKlD
nnFbBAWD2q6LreKdOBvSVVxNfQGbbBpb3MJjdqaWHciJhxBoUCHOVnCtyGlhEnqL
VtcYn6fGnS0MGqqFTvswE19ylo39Aas7n3AzyxZTDF3JcYMI8OdQczKtTCBQF3C9
wBgg1EK+GpJRoy2HwJJojgPyvJktvGJSLL5AzRkNXQL2ngtFYgBFyuHVTCdoyZcx
Hw0vNE32M0x+J8SeKivMH7VvG9KP3mJyX/wCREbjT8DAHYZSeegPUXLqC57K3VE/
C07lWj2gV40accy08OZEti1nxCOZSYogbgL4n0B40wcvCR22oqMU5pxFSFK9yOk8
vRJwe/IuZooYwHSUqwBeXi90+epE5vYmoqkyh1gxbBnsYiSyJmBg1QjDHrCskilx
xsFnUajRLb1u130NGmXMWd3SVuY2CLZUze28rFnVjhN5hJTDFnXFmyYTdHPXEckp
6t06L4M02edq3eKY/7q+4K546GkiB+9Pgw3WoIbGGkjLfJoAmjgpQVjvh1801C4k
xDD3fl8SeAhFgQU0OWEaCJD0+Kdglm9Dh5ueZ9W9lIc4fOCTVO6IGud7bOBd8c1+
pfyozuGInqWymKHKoF/5cbrCvg0MnNfiD48YGhPYYZ1yWYnOM+IXOf7WmjBDZcsa
Y7fkakMKX2PmLgzb+0cwfOaWZYZLVa1YM/sIvnwGOVsYuIuxnrvXb+cN9ND3eQIB
90MmiLUYorNmOliTnDpAN+mrm1OfYPK4zeGAofSla6Z/S5zbLSFMxWF3xpZpE/Tb
N43Fc931Vw9BjvHJ6Zl6TX0o7RtyADZsjHoJfKp61/LoFngHM7o8n5vdNtvrPD2q
zqPOfbtUl1ppj63awOvOW3Y+D+TQ1esNl3Pvr9x9pODCuoe/DKAnmvVoUJoIPOJU
TJGjpIavnKfH2+V5AaK+jL2uQ4/a1Pw9zDVg9tMF2SoS4qBfvIlVRHhKYzTJ2y68
V4pKHS8umY11rlMbPcfeiVNbg5rGMy0Bq8ndJnwk6LuWpg2JWcQ1ZZlGj8pRRUfg
aUhVfDapr+28pOzEtOLoTJd9XdQjTgETIC5qAHyIkxgraYrBhI61YCIsd5yNKkx2
VUCxh6Nu9Mj7ZFC2qXUBc3Lo9Oonl+fp4uyohESh/XJFZ0EevhetriYqTBIWLWeH
SRGZ2+V5Adoso3hHv+nIREtDo7DO5D9OZ2ZOBkQiTp7iaIc7xC4mFgcl4jm5eEqe
jZpdriyp+pCWRRMt3YqiV+qdI+GuifjQVlgp+3QLyT83yoyTUyW8uCAGhZ/8nHYV
/cREC1Qc6v45L/ymleAOcKHLxmTzUMpfBYnANP/j41m8V7I+NgED0x1LXX6UyQif
T/lvCaao/Sn4BIWwfQGvbkJFgjkEnOscWvjq+wva69LNvgquGx+Sh+iU10Z+/9iR
F1nZxu0UsBts+Uxa0aiFSbxpdq25nVm6DsEYEJJ/0+RWC6VVhQqiPEOgMo0C+IZX
nozMbRmvHPEzwJZ4F5KU8ENsgLJqUC7T4s1U6r73Tw8ru24ReZkUw9GdmAceVX0Z
FC6E6VVDG0Xvz7PY4Suzs5lGar0BRj3dmp3JQFygoO9tx5fzENVeQB7DjVsF+fZw
WfEtcZ5HgK0vVnkJt7Rzbs9/H5ami8Ftx66pNgsgIEYlN5eUJUWSUyKYlSv41+77
M2eST9Zb+b7uXX7r52FinShGf10/Aty7jN8adOopGatzYSb+v0eA6Tcij0QghZDD
kp2e9fbprSiV9k+RKxSnIZ9HWERQid65ZCDbDyp0YA26vNr6pUUYyy4CMq7vt3yu
kGkr5Lm9FX/2J/cin1QNWbVDDfqn0pf9jjdpw+NZWK7mv+meYxNXl4pQW1/0QyU/
M/Vs/Ca0PI47ZyXy9mFoq9hvdpA8xPAi1euU6lWeUojT+eMAa1rZMR2rRGlr0009
Zb/G5JCD9uXgvzCBb7MDY5R/mHQanUx3Q4vAYsowIB5x4o8ndQSvOQdYocco2Mcx
I3Pwk+PZupz3n+RhoqkB3AIswenJurPi1vrZEe0/oUDyJsZ23zfx4avx91FReCh/
ckWym9hhnGLTN8jvRE8ZcXaOh1j/2o67bAw3I6XSxpXkLwuRgjNzbE3PjmhQDphd
BS3mIyLoBzI2GsTnOGnjcLFtZxqh79/6poe7JzMoiI+ClRVbUez+zKuVMYGgTO29
Gs0RWJLrE4mka1alxQ/sIF63cRg3+zmkGD8m9TO8mw3WeZkJURzeYQjhl3XJTOkB
YQqSOmNY6FocdZWApBtDJdYUqbWP3DZ/7VIEJRDmNdUb5r6KrZgn1MKtE9EFshzp
5tsoT+zGnpVsvkHcabInDnxQjpOMClbR4/nCQEqxT0c146zFaIsDC9jY1+8/AoyK
/ZViN/yEqq4ZmurXdWaQTr6be6LX+CYyhizfaqeP4A0uoqKgPrVcBkP5tftCMrnc
pXkoaM0uHGDaF8lxJ7r5cPT0xa9yQ3F5p+u30kuVrMeaQCQ7+NIaHW8y9/pknT9x
XKWCH7CZoeEqFFHwjN1bH9hgxbXnBON51bMWxp4RluIzQbNCLxUk7DFlH3osDLur
GvRR1l67TRHSaBi1RcjA+d4SfVjOhEFCSnvmHrbHWnEH0IoFg5cR+gT1HC3gN5hT
qpwBZnm8n/iwjQhO1yMwXsQYTY5aswpwZVoW8XvrtCkjcEl792DapSYOeacWiEj1
dMVlTrM/LPDR0GZUuMYnxiLygQkD0nUPCJ0nzLq7zLzTdUb1haGc44p1tLDZimTf
+goIgorSQisQ3Qt798vwbB7nqBrGJpcjsL1Q1xy+5iARmQfaToLZPQXtcxz+zzLV
rHYlug9ckIUipaJciY5ugc5JGiZq0s1YlrsdjT7XSgZu8fCsjgPeUHU06NfvCsmh
aj8jotPA1kl/BKIfzcrI9ljZNZi+IAdOI6rsg1X5I6+99PUkJV6Y9QGdOHomg/Nm
G1fpV1EYjzSy/F8F9N7MzoaC1ykYfCwmbVjS2HkuHpwuRaO2YWTe02hxz4OejPWY
IJr1bfpfUtkRpK+X6fWrTR55ijdzllNGSy1iATNWTqINDP+qnB1HWbPERFy63Kxo
F1p7cqKsPP/URxmS8Fa2qfjtRA0KzjXyQe+gTxY15KAteNN62hxfmf/oCzOQB77T
8TfVMkjVLLrh9l6g5MQlZXwr/2BCHai/ZUZHpqWz/4xKOj2AzfM2tYgbdHARb7IW
7Z5z8YT3i/bPYgI54A3/T5iVmOlmLsn68UJrzSJuRDp9fkg0YBCiMqMOkRfXi+nI
Ybo7mkBiW5L2u9qfQS3Yl8YtGQsQzkb/emGz7lzE9pSu60ty1hDymdlZp9RpN8wE
I1NtpHUqymWIkVm0P0ChQIeBXiV7UM92ekmr8aSxy7oyisRs/wOK7lFjRZgtVpyG
8y158gaQFT5DZf5TBwWE6kQcbARThAvRB6ycqRf1gssXbJFdmys7KpZ7AiB/2SFf
pJO3AZmToUWrB2J4Em+H0OO3Z107djprJB5Sk6HsmAPIHr4Zy3QopBepIF+B27eh
XHO2LJFO06u1R5oi9jFwYgqZcBmnse/aFrr4Odk5mg/bYe5iKa/nRvMLUBjpyWke
HJ+7PS+TjvQiMpfyfOOkRZoGceoGSzRnOxJzVkg5VLZYqcsHHm1A4bPWXSzlNrMe
uJslrpX+pPpaZc8L06T6aDq8ARrPlsIb9QLQzkeaGT+UDztDbcxxfyF+RE3KL+Bl
wOLkvcOUGrMlqBVQPwEJDAecYZAx4kTjB6899MWDezbN/E/GUL5bGdvzp7jlYozw
r+aPoNDHzIvn/l3xvIXdaDLE9R/SbGzxqT4bSFz598EmJzShI0FHSzTL7RQvkbeZ
U3Gc5AJx7nd0ePI2vw3IMs1xTwI/po4anmFzhes2k16oJXoazrI+M59cQ5Avgyny
xrqEpda5KqH0ERlWSHTjQOngpii7rkw+rtFM86rMuO6P2YHeFDoe1n1lLjcaUUUV
ucQHpPQNSDFaBfWQfF1WVBpA1HTHt/vYj5+x2XiXSBO/0Sj4JEBf8kbh2C0IntHT
uoWYtrz9XpcneOZ5h79kRlXr9jVI0jqM7iDHVCcV6Yb6SqHOolMDPiva56z2tkYn
8DdppOwdVcMgj46hRmDFaWK7CSCJD7IKUDApvTRTSDXehdXHjSYHShnpjaWPFK9F
Zf9Ns9TGSqEQOxxtSnO20ZNsDnUFudWcCtutxRjIkjfVaeKh6X8d04UGn4FQsCPK
e5P+7KrOiaSBBsKxZmWMMsrbDpWn7cCOkDhxZBtwIsB12zlr5R1Jh9weY4znLag5
wu9wg8/ZRKqCLwFre4Oh2KHB3ZaWwVfcVkqrq83w9SslnT0ubU5xQAxTtcjGY28H
k7V4jJ9QbllKkXtJTdlTYZz95rSNKulKutjPm53dQMF4jlmJbdxWOMcyQo1ftCUm
1L7iLBWSIRZEZ8s0d16xDrkrfqsuYsybSeMBimUKYN6LWWLXM2cWDaRjSlLjPwM9
tdSkni/76yVR56zsUKs/tdoyw1m8/JHOIIjIy5bXCvcH+oEuXs5SpZvoKewRGKT7
3t2wW20Bkf/sdjf9VTyEpmZCN+lG+aRoi4mfg+imQR+ENxfPPQfabVuTX6qNBjRL
Avz5VpfSfJ8N4csOgHMFhCgGx2T8T+AghQ/Z1ohukXMbQUg+vL5VHBaNvHKyYgwS
BF/W/Eklfrhb1QJxPZg6MJn61906FFawvB9mfrv0SxadofhOkCvg0+eE4EzznzeN
LNkHVi4zmD2XyUd1Y0wAhvMKo0u0zJxFFk5sUQ+dlUrSo3mpnCmPh5Ri3Ur1SMeQ
ofbuDiLnqeyxcqt2fJRDAqHghoGBd7CA5xxlF3W77xcuRUvUjsbsnf4XRvyIcymT
hb7zGK9l4mp7C9FjDjX/HLXQoYVUSVaVq+ah3UfxPGbp6hfmAsC7RgXsnHtctnHp
vD/f647vuqOZmvSwvBn0FDZ5MWm6mNH7V88DyJi8DijQb8bVsZCp0+eKE5e+Ng3O
NA0Tzw7Iy1eEwxD36x4VjUQhksfJvLut6ROVSohEU9M0/76gWXSRReduN8qfhlKm
3D15OY4pK2RUdkfubX87gH+1EQrLG054iZ4d0YkdRjlrK2co8TZGtTkbK01CoLTz
jON1EyzYDAUDWrRMVb5KUuM/1yJVeMHQ0CAdq98xZkj98qXbCACR7fl/40dkwF0k
5JUlmIdcYcmsFw+lkw5nds8IKuers5S90fO8+nsliC5GuCok3ElIobrAyYN4zzOa
RVFrbmiKbBa5N9R/x8c1pYxFOsTNGlvxuld2bdQjEx6wXwQaV/5Q54toszqth6r5
LPQd61qPgoLKRxn+qzciQIHtKXC7+9V2dM0VqTMgkFf9uFSYilquKy+qee7fhja0
6uf8t/G2bwD6UjTZVap4OuAWyL2nN/MB234mVg1gNIV/ZTS0sggE3Kgo2SpL2QiZ
zbL4GjihtbsVtZ/NtuFy/EIR88hSb9T7fSaAnnSESVp4bGjK5KnBk6QzYMbs1oOz
nB2TxZ+0K2xfC5RwFU5sLneKesX0lyV4nLZJsJfuR4gHWbqcHgcXuPyZqzPQjt0a
egigth1dl/mGrS2741Ix5TdCVeZ6V5F9Z1HRXzG1cW1wDdxy3FlIOyzKtMdU+nTS
g7vj5QfGwuVLemZgAK+M7O/jmn7M5Yey9gjGAKOaxDBJZTIdDI0vXAuOmm2EkBiW
YC8dXpUY82Xurnsgx4uQOdLfbzmqFoQXwl94TgDF0/cJ5bQ87hkZOObpn/QRXatD
A0ntrOV6P34cve+SLC/NsZUQpudcI791Jg2Y4GF3zMd5UKFdGS9GV4dY04ZJLfNc
OWlkK3bIS1Ku2yYCQ56oi8VRmIKpsXO6la4lxBIlB5UI44+unmCOT2TYWMSEG83u
dvBLhWRXMI4HtcoBDwycgrKaVEhOE9O3vXU8kpUbALELbdN2ECdSyrkXTkdUp5GF
oxOzUkMNssLeEiC32ARNiQ71PcDHTjA3YL4KJ1sxKe6pstoxI8EmgrS544OrXvHQ
QwkwWstPbX75QhIBNt1Jaxvn3RbSeFYI/7K0qPz5k5/RHNthYWmvFEeXfnZzlzTp
lPgAgJGRTvCw38WjPemZcRQ08dJKZP+kAVFz1bn6Sl0DbOX/jsXGNSfuYDL5JYvz
bmWcYSGN/lCO2ylw4b9JBkTE72p4dGONiP/rFhFJVjSN6mL0dN9yPfyqL39xlwdJ
wJ+1oHJQv6iFugJBZRkwnobju2d9RUgLSFZTZKjV8oobHcjh7cnPYkLQf5K01vEi
rWvR9sJrWJAwWh9WRl35/lroirunu1k3QQRtVgZHcu/5y5/UxW9YDARiW7dxxZxN
eeCdlETjlH/kGSU5gzowPcLIAvhGLdLFqRl0pZt49iKd/2FM2Ks0zKN1HRgkJTfC
gkRHOIA7bcUN5eVUOfFA9sPhGN9jvnTpreZO1q/tdkm/a0swd5EK7k9Y5b9nq5t1
F5/62rU1FjB6xHN1ZuCzAoCP8M1Sh6Y4td1SvTVBOpXkD9terLTWYcOrE2SG8uEC
pFN7QmT2666NluyZcdLLtAHgOpSl0PtoDAfbZarZ0DVKxjiEfaKuvtRIysVFHjtG
cRi2bqvmNXWwpllmPSq3j86gUm2MB3+fQz8eo4QURAdc2SATrVB3H3J360alm5u+
r0pqxxePDc/I8vEZuVyR1WLI/yGuHFr8NveV8OZrykjpPpMga4z+NszDh3/zYDtq
C8YFuIhLWB/FRsi3XMwHyWUuYfSyMG81O9xUzBODwviuVpT3FUczIiqnNT5+ijju
jETc9xuhfWXRCdvqnW820/ta21mzwe/nIu8rBsuGi3rVTAlMlgKFShSfUXXhsyUV
zAyyy3aZZ3iU0L+mwJAIZic2G8ytT8XPtHS3s0csXpXZelzFSF/exsewm1wH4vtv
rlVraFL99JHnoepQ+MNPYXhbO7DNi6ESoN04LXIPxu4PDTYN7l7cI9rzQQKEatSw
m3v0MH24R14jl/GJXJJnAYMyyyN8zMZ9yCnn2ZBn5bc1giX8ugqdBwMa0LFpoq9h
nEmztbwQXHxEihUnFH2xbKd14R7ubEsVcVAttATlX7+DyiyB/hfiZUjmAaeP5M3L
sexxCUvjXRlLu9HdSAMSoGq5Whk5qqCnE4glnYCB5zCdE9c2GGCGIv4qE5rA14oz
rCBcZkxeMhivXlp99AThxViGQwhNdFK38ek05tl/4pvEAgqthBWKLwZckZKskYhH
QpKzDneG8sd3GpuiyZdiWT07zp3PNuFCdna02kk7GWJ8Pni2byYFCmjbeqGSkW2T
yMC407pvWKRN/LdvEa6Jtoh0COBMoy9hkbF3Ua2jmWo6OdtJLZUpEgl3dtwlMluT
sn1McudSPpDIzMm+Ea2PaNZyfn1wD2wFQDyyrRrI3wdLe+OEPfb6FWzcJw4OWeCy
wruSvWBn2Ok/PglswMPaYhIHdlx8+pbOw0i3fUhzIeQ2be9Q43WIGd+Z3inrf6H8
Oy6ySwJuKZG2Dp2NQQ1eQxW5IXqnbOVDsGcniYFi6YKUFtWF7MvIu/sVO9I28ffK
9hAYOw/AZP38TS9PfE0liqibjOgIPw8FBpPLL04LhkJB7qheP6ugY39LNzDFUqde
tr8a2QwRtPDosInUT6ycosKldyyctCOEFNP5iB3Cu6iYmjiwPVkwsSToKvOUkePI
hXmjqoKLgM6G9WuYvoXMn7LZB9OMRXmWyo75pqpBzFT9L2PWKF9bSJDdMI4Uo7aM
T09rTCFwVvx+7MrrPe1kis7/sBaSuar44/coC6c7FKiFXvaX7i0aQcAjBZh/pJ1Z
z5u0TZzz1UBL8mjRT7pR/H8OX3iz3Kz2/PgeheLIbQzr5vbTU4KHrWjx87CFEu59
3isbKMVbF2YJqFdHED0oVdd+Y46OYLyXYAY4gGp/RXzK9ozdXArWpUfe3qof+zmm
hZMi4k233N4fpzr2vm/qDaHnNyvW4tgfX5dbz35g4WWukxcgIEzog2nt/Llj2JPT
8k5BmPBaezDaSqmboBxWy5aiJ4/bIal5Uu4Jxw0FR2OMOuwRSV+/BdaLtMr7Vt08
YT0X3EEBKXjjurSdvbJNENa/61ASTQuFsCrPMcgPaekJh6Mij8+bgC83Ey3CoRRH
RM47Yd3DSDc7xw/1RUIV6rknGpAfgg4Wp+N08sf7AVsYJ0rkkEj9bOC2/qckSS38
MIw9dkAcYChT89vKMt+XTc+kQbK9KoZQqk/+svK9scEyC/VZ6szmMwzzs/Twkb12
4GyFAg6ov1dYu3Y7Y9YignTa+7/NamYQ57R10y++bJ9g43AAWP4fooFcEIHWpmBV
kT82ygszhomkXutwOzy2d0kKCyfcPTebViVeCSe1592xuAtrdiKp7TrcoEbHBD0X
wcEZ1ueZdd8Fd8+40x/wElh5yDoeoHSX6y4UCLXfxwl+hFCy8ks4nMhqu9CHiLIP
DyUb4P6pK14eVeSqQxt5j83YTEBK5mBkqGx+ksLOJ99kszbagr/+D5j9eq4YG43D
XD99paWQjG6p/m13ABww4kjalI5uXlmVRCLVNlmqxKV+65O0aTkZ659PZtSRSUoq
k3pxnpSFkvtAICR5yMXtHltJymdWlhZz0Zvm5NfsdVSiVdJuTSThKAmkvqVnaFc8
EIL7VHExnP0oiUgt7++FPaLioukfeC9BVMiuxDUJtIHobvo89hVtBkevQsFCFhFf
SoSN3hlTwldgzW2VsG3d7EG9/7ze3Mtp1XRcR9nvcpjoKkvuBNTlvgUdw/PuESql
EGtXeVH3M8FoBIJL4RJQsFCpxmSus/fJSZVFHoO1Fr5nBRT4BFC/TXCNkJaztCOT
w8dtHAlO+4bOU1QxT6a7A43udNYhpRbmhEfR5sveWgKBYnU+TkCyb1hpfRU9iA1c
AEKUBRmK5GQyzJk9wDWbu56f1Y6Aqy/xIjesYquRWjhT6zwMhSkwGDB8NDSe3NFK
o2K67hxtp2+o4RUyy0jMY9J8xmTHAYHhv7TCrf9Sq2u9Znm3A3dEp76c0nQOxYcQ
2MzybL1R/K1uqEtG+CWj0Xv0Pxl+0pvuXSp6QkhzBbm+tDhYzpLGwJSlKCTcz6Wr
0O/mJG4TQ8L5ArWqeL3u1uWprSLO+uF9urW39i5rBo/0rNe8uH7Q5Dy3fkS0UaAa
D0khTqGypNsP9XaHB0IH2P0hJ6R2o/O8R+RKTzHMz1RrmV/yBlJYpJomRbzH34cx
tPmYrSfQ7VZd8YsaH+zINEK6056OJeosni0ZbRwrx5TqJERJWtGT7dP8pklUmOuO
+SF/zfH0qfZtJd1jM8UXV5me9MN+TOhRDumjUGZIj/vDpYOExF+8A+hlgkVnHJUQ
k8BCjEk6lkLjeULQeCMlh0BO8Bjsdz4h8A4C+vKbI/z2Hwhv/oLl72TclbpCSVLY
LMsnvEVnJ0QB4KaUFuAz4IOSPAAb4IPChmZVZnEuUZ3eg6qypS2L4aOvYkbyz9OQ
RP7ez0TjbdNDjcZpNLzDdzw7tr+hWNnfBGXsY6WYFq5yIuRHOWON793rAhXd0ED0
tA0efzOXLaICMZZSfKWItKce8u9hOv8aic+KKSWLjbtiiTAU/ncbbj5hmdgGKh3N
X9HImXSfKLPUnrHc3e1kPbK/dZ8H6l80tYdjzMFSC35AJmuUIORulWr639LAw6qL
6N84zECRntNn3jYlJ07Jn8bNezLoo/g7c4WW1E1/QKM902YBE1qT44wk8m3zLQn8
C4mEjF0cKcFm8AyuiNLQiQBKAUbWCRSAXRN1utnJapH5sb1hg76616AWVyGu+T5y
xCHT3QTUQTbMpyogkxJCxxbGNZ9I2C+d0Vx9bPx+5vrrJuH+69KM/Uhh+XT+ewx9
Pz4wMmzF+idQ3zK4ks3ItNDD0uQ9Li8clv9ANbm2VT5sQxE0jM1aAnsFyFPveM4F
R8Qs+/0KSrihukurBGTatqNL9v/DdO0yloNHn42v0JAiEw/X5CuEng1d7MDhWMYe
FDa3d8qJcSOkDzCC7SFQl1J0hChF3hgx9KgLJGPVXNLn3/GF6GjSxZG6UqnzvTTN
lJAB2NjuaeCiZiCJrgTwLQ9KHJEwkuYn+x9xQJ/k7Jx8YsKQLGncgmZT+4lJQK+D
0sayzQaO9eatXGTr7kBjWG/SnD/8984s8DKkyEkwTr/4aYqo38jOCsIR1f21IPE7
egvKeooERC23wnXZUizgNkSteW3iEfHTAtHvZ3DW297T8WwNfZBD6uqlYwpvQOzQ
lZQftGt/Wz6CYYuCvQXm84r6mLPTWdxcfLnp+eLuxhtUZu8xwCDRB5Yk/aznBD4K
BEEQqoevaq+nqMUp8zy589Xv/Y1DosGc1tKxdxR8dFL+l5BYb85TxWGPjSSInYM/
XUe9YnizCPr//EZtAHIxHeW28JIoHevbQ2h3TksOzLdsW3gPN3IrrDz9VILUPVcJ
KRf+N0Qp8B6Vai6/xVa/989aeBZTW4aNRlUiWGHSfQwUFdvXVcHDzb4jGwtadTfm
QZdgVeGZPMDV5JoR4qZXyirmLbKKyIJjlhvCSOZxS63ebl4w9+V7E8y8c72rzpIy
suvpHQO+GrXWPr2T3Zm1PdNMYeaARkcMxcklgqOrbHqojqyK6GtdnSCXDwKkRJuL
etS7YkOyBb7/pzDhH5ntaOlmfk9VI9q6vLw8JQH5erCwRaemx7e2ebd8ob1Ax56u
UkdmZwOZEX1QQ6IKnx+lL9wTFTFmxUADCK7uHYxMh19Voss7SJUofXoaAOz/FwWm
VMOay3txy7Ss7RPnxRJkmMF6z2/6Pm8NQaYzqFpueafEp952hBBsfVsq6QngiiAf
sMc11/j+6aovVBnfZ1x508b8gbesZjZE7wvgOcDLBr+A8ZfXT5LhddcHFKfSulNR
rMxQQi9Wb6Nhh+fLDce2FaYHTZEe2Zhrmk7kNpLABx+jspnBJzW3WXFpShdIanB/
Qi1OwWyXzO1yJRKAE/GxNsmx1qJ0X12sZYzRuAzSCaV3f/WqrpmHOBw8DkgjSPfg
+3q4/VNmdeaXzOmpuiIFEdg4gmyrht7cj+NHTVO8X/lEqwaJJHq1Hin+r841DrOJ
okzeaZ+mDMz4MYZqNw/k9DIp2k4xsMdO/aKOxQVWvd9z7nnAq1Y0vatksG9ok08W
1SbYfSKn5aCsXPTm3nE0iGwc3hsYj5rC1y5tNwW37vXb7z9SrfmJ6v1QC24RPOls
WdxQgiGNP6rxHjWBFHQtBN1fF27rz0OQDXBYMbILwRNLsuEzMADRil3/GYNxyxeW
H3SvbTuYlUc6rz9OtINDHoHLgbh+H04mNm9H1O1YRep+bYrhfjnotJmylVZLA4gX
L8cFyW6BCM1R7xHXuL4p1USZfjE6KfS1k2HgEHl4jqfGunC5USmMgBg1dM8nYu7w
epeO35vYTWuM1hpPTmiAtpYXnwiYwIIKOe1nCs7b29F9fHNWTo2mgh4iybMN47iP
PjtxtOWqugUp6NoGcMAK8ZTAXelTNZ0GPCGTUxP8Uznwq4wGUcsp1HAqB0K79VuN
dpVttMtkBZMh7aEBxexm/ZwEA7op9TXOfGgOxGoCJmbc5fWKlbhXH4B0hYNtGNq3
/P2yA4759MwwOUj0INrW/KH7CqdDNQbunrDbL0dODFbmLBQEmYJ8I6va3vXcpAGe
VVbIygYPX1kEtJ//UCbapvEVayvMFFPShzSO2Mr91FIqFOR/ZRpx27nedqFN+ar8
C8XWUtwNgHBevgvkAa1XTHCcFHxtrjZjGOqXJcE24MyLbuVAgaLUF4km7IMlIQjj
fupgnDIpUUtQjJ2d3KL4b0djrV1KktyXNd6CZS42ijKeOVAal8wIDEGxpRkFaNoy
2Lt9Z+C1ffCppU6hMaLnaqMOtPyOiToP/vDOqvc2x6CWCeP6iDYHkK027/0Vzioc
hR03I5+Kq8NDjLgKJAq3jHZuPQQaKl0Psw538Dvn+xYeasopxXH6yKCfXDZhkfuH
euTjDjj79UNJpG5qKgk8+XKR9dwA3rt0YyaVpyonMbMwFPDXQwUuWGkXfDnq7+wC
iEo8GOmHEYwqE/bQevfwZBgacOCrqRplKUDIeQgSkoHurGJPNk+TEGKdceLkE8Ed
//19CAcUVayIhQT6gQjGbLgYAQCOm2Ndl8d7Dml3kcVK3B3xsXZ+tpTAVLDPju6u
PIUraQPUUzRQHCz7kLr+d3OwsWk/LqwuZJ/GCQkuN0UXD4/4ydLbhrQD7F+Ev0hr
vMBjnZBX6RiGcc3OfADUqAfauA8l39Y1n4Dkql0yrTNiRVZwqq4WiNYXKAvyceI3
+piTHdXvLduwWmOzJIerTHod3wH2o674HlMX40XIx7Pw7HlQ6Rz8tN2OH4YXpl81
Bd7vHbyxN1bX+h2wh+DleRohMnk5fuGEadf8hDigPWG6ho9/2NTJSS0zdh2XDhIs
c7aBhHFed1CtyctMR+OMLPwzFzzHKJmBTtxW4A7zyGtiqf4/6tLx5Ud0aUp6MkNg
Ka2bIeiIKOBgPvFIRirJrRnURQzkgzR5Zmi6iMHpLEBHoULD5atMhPvk/ErwT39v
L/RMPtXliCpgwsrNiSaNghGQBKiLbwUJGsKl6tPruecQJN/KpovXTZsSzlKUZWxV
IqjTQtiVt4l4zEG47i9X8ljR02v/DhI8RoRgLkyBqJmDsVvdlS6Yf6ZY/hV44T2E
fNo85/8MVZN70MBPQRzcyF/LGnrKTvibPWwBNhAOrWs31JOsJERiYUiW65aU+9Nf
B5Rm4Y/Mdq63paVbq+a8I+0z9snBLB//WDj5SV12FgJbEyYYFm/v2NqrTN8S+Ds0
ONiCM+qos/REoiijReXDiFauUOB4l104PBi90HaVyL16s/NMHtFQqRr8OFJW6Pfl
cHhbOQBIXl5EfbbcDQQ0gwR39+CMy5nyeW1c6JGtOuqDUVnA0LRa7RUxEdcnHeT8
eJH3ScADw32tGb9KsHBBsKSEiNrLbxfCy/RDPMuT19KU1lOvZJhqkiONOz5dB9j2
zmlhuUNddpLRT0CYLsol3r8AWL5ioLdlbjJNeJhBwbYNtdnIvexPA2ScmDXoVubc
pXXHcEFLXPIRQGji2dDbDPYmUXMlIHKZyfPiVnKNyiCYtnUjLFDE2SRCiDk57PBl
RAvrD6G5kNqSfrswvbIqq0Xo9ANB3ei02OSZe5labKx/ImcPXiVCBw0vpRzgOxt9
imaYzgM8bw0SFLH5X03QHJ9H6qBTBH7d0bMUv3PrYUcZ3LjTrB0Xi/KGCD6L6AuK
LuZwsKww1eA/4GsrzXhZQcx/0NVi+tO2R7zJu1cyCT/t0qrTxq/w0B+ETc/h/XQj
o/Emrwo04/V+UfD8Qfv+vy3pp0M4/kPs0HQckjc5sRabxXNQoDM3Pks0f3hWesEs
SAJE1JEvbqYv+J+oXXK5TnJCpX8F45XpzW2aT9tae/oS1TgXIPpOJxwnd5LHG3qI
cp16er7diBzp+4nxz18pZXPL56C0hwlN/dZLPpSXXdlSLOSbEv17eCBqxLYWWp7p
rD8YFzZNkD3dfhfSgFyttpiSxjfhv7ggimJ07CjlCUwjOSqKNn1wT1RFPskeCLi1
1rLyN32dRtFCEphdMARrAqaVpvmRnxAWa9QMxc/gi44nr38s2ShfnKsR8X47ex4y
RFNiVcpuMk8GKueKW+R51YUj5/Fkc7BQ91bO56rag6+gNKhMr/NdqVZjPim55moJ
TjRS4WAIyhoEvXlYpf1Fx6bQwT8MbbZedQYl7n5NWhTuo1VkQRC+untlwGfsBpoc
VD2iS0ojXw8Np8h5Dkx0PxxAfmuHfM45pWnwko+nsyAFA6IH+H2G9NFAvrVWaD1b
f3C6cNKoM4mmiM6W6smYiAYCBgMBRNoFTze9uHn0oNFyAdtndEzUHKDlHlj1aY1j
TriW2f0OEt7+HBTEH+KOXKoFg9s5rV8l9caSXrWJwnOgoU55HhlBPQHpP5xM76md
jAyXjd7mKbNlu3dho7PW8ply2Dus9r1fYhMjqOctiO69s+UZtA67ZBS6LoF8SmhQ
Y14zur33y7iC/q4pmrIe4cawLGD/P01BFJJvbHp492pC9nvNapYoAAjG2GPjfyGb
fsQ18oVfri2x7/PdtdZ/7R0UiqihjCK+TvL1gmYo3nYI/1YnLa2RSWIdwfom8+jD
/vJkkrm8TV9Og6gZtkxN0z9qvks8InaDaR92mL2F+xta2PBBMjXUZvluHxvXm/HA
cQz+vYLg/ms0NOzlcXgXakg137n0atT2SeRB6V+lx0iS1+CdG+khsX60n86Jfn+X
/XdmhP5OoE4FljlSQetRweCaMxCwPcgFV6JMaQHt2NCE9ZB9nlZlIPCWJlFmj8zE
T+BH+AQwNWdTngHtUd8VJ0i28yEzhxYyogtzVGquV3HERMrAEGKz6PcQi+BONyff
3trmv9uoK0YAHi2NGBlz3Hr+XH6d8xGX4L5OlSP21tECRmx4NXj3uvGpoXKIt60z
XCPA0pxCovDbgXvKJkxalhJJuPwYzcY59aDZM72yI0fckPJbiuO28Y70JtHwl9ZW
2ufbdL/DSFM39GdsdNQDai23AWfp0WYnhLTghJlu9FLxyTaialPmne/KSYUeVaOB
tFJOabLUMGhvyqE38dtqsSjsnXSSSQMDdRiS/l2LeSuFpWGo7Dyb0p/FanKB8NnR
rVrch1hHgBdVi4iHDIqqviMtVxCiQx6Y/lTKs2Fa0SEdL5iA2/byX5e6RrL2MefF
prxQUHpyxQVdHyzBA1PLfW7OSYdpLA4y5APklMCLyw7lIk6o207RnmbpzWP8v5Cy
cIRBemba9m7aNsH96sTpKCfcr1SOacjhbUzrLJcoI2wGzT16bBxcQb32Z9Jd7eiM
bQrq3m9m2Ll1Ox14VTcdpy2t1E/2LoaUd9Qi0Fi7AZ5n9t1hUd2skDdBZbynJv63
DUn252K18hk8j4CoDMNRFC7GWq4FCWQ+UvXyaf8T3lyU2YoIhOX8MyDqV/gs18vQ
HjuXW1jaDYGAXlKDau09yvl29MHnOe1dOoI5MSRDTBP3AbxazKvAnJ1LCmkCwanZ
TYVJVLYxkcuORnzZQJcn2+Kzc6wbAAQqlwfPyNzgK0cdjuaiDun3sgQkfjGQV64M
tClM+totB/htHo5/O7zqgYZjpiLIhiUSXVoZsqVaBvQ93HwPW+oXbTtKsUkuRYvK
7MX/ZWEhNG8JoJ4h+grliSPt2HEiLbuIgg5baWvRkFgFq8sQlo+NjaAZGVrvGyBf
m32fKr+4CouokG5AEf5EjmLX5IapbN6ENtlBu5mQjB3GxihMEOuh0MyiTKCHXV8H
FOC0FwUiT+HS/F5mbopA/mKHJ7SAWds9VGNWFqFJkcWYzlKZKVyu+ADjBMk+M8w5
grDvV2UkVOTsHneIXLWILDjLNwMG0nZrr9glJwc4ueRvg5SBLVkz0GMRT/kKkVl/
0LMwxKLGmdK3Q46KDQ3tQq+iUXZJ0wUPyJyvxD0YSDfp+OWOjsiCIi5BKDgZOuGe
+cZ1/96V8esP0L2do9o9O7FLyxj4LF5OG5abwMtu3OqeRk3djFCfU8cOLUchuzKu
ofXKR+fI/mUfogxwYU5Sx95rdk+/J94n1D9CDi2GcxNpMg8RZN20TPNYx3BrWkFB
Zghl/IuEo74ddEtBHe+tXq18gh+4wD4HMY29CUhH55txytDf2xT1sZV0d83BIyVT
rHOioMB6r1zzowTk/B/sX7XmkgFc2N9aTyBqpOTgD/sD3wG0nzue0II6jPWmSYb6
dl3HqTMmCSY+r+iGzu3oGG5OCFxpXqtPnW2iZtVJd8uEo4KBXaQWQQa3ApWhrjlN
UzMfHVmd7DCZ+BWdPl2EtbmI3Pg28db7KsNY/Rh5TAu1H2UjscQAu4Wtug2SzEjy
FPAEnsnMQfBlOtr/zMGDJ6VNeTaqJUyYlFPQQHFEzotD22NprCuLYI0ON9ZtC2Iw
alboJfBojHuKD/0sQlwKS0kbNZS3U17wb7OVqyHWZuFOsnt1/FbIe5JuVc0nSju6
i+R4G3yrt0gDtLHIj4BmILAz0gC85FSminhQXlDpCGMMuf8jZHkAhFEi47f6RE6v
tyyKZkFhHkPmz7z+xbupCigBm9pC4wjWv5RdFWDoWHuVm0rqUvnfWJsm0tgzQzhJ
oOAKxq9WISoLcb8KnqHrAleK2z3PWDEfdjRCAzzQ3nrSRNbDx7WzirOAX2Irzjpz
Jsiw+D03zGp2ibD3wb/BhaVHpW+mbO9m2lvy71zWR99iXJoK0ktMH1HWbGV38jEf
jKs26sBP8AI52bPO8vhZ2AibrF8BcCHTVgX+TG6UBmFp82AFrbfJgNOYck30F2mS
lvzIlyV/TY9GbacaYei9lP9Z1E46G41raBXEzOxN5tFxHhKfCwLiOHPUtmEfNwg/
W+GZh2rY0YfeogTI6GWz+HpGiB2n/HSoMZAM2l1Fb49dMgcxJ4s3nhhsp5/cLK8N
E7EihXSTZjR21ZOZ4PRanQuGVlECAqSk2+v7/FgRFlgPqLQCmfn/c7ZYYFTTpTmU
1egsF8gA5bohKW7cKLPNjwcGRsbOBakNRvfVod/tIFXc9JVj78rX5jM7F1emYr7N
dd1KPdJtIKAOGmGs5nWz2dMbRXvzLFS5v3J2PAjs0TlInuR+24CxLCY34deNi2Xj
uWU5+MwSX9SELSq/R6j7GbjRUDPC0s+eRzFlq9Jkw2JEY048as0eU5SryrfUBf+q
FZLlFNHQxRe70rotvl1MRJ2W5P4Bjbiil2aAbNoK9m2FwxYEJegDClr8IcQ2fzAF
tEbOknkw+BoQWR4hBMOHpE2mC6m0L1ktLxYSeBLfg2IJnziaZoMI6xE7SR1cWRU8
Z86ryVBHBMfGq84f5u9dZcvoPweG8lVKnfNUX0F6623dOwVPbFSVPW8QcRiXvYKY
6u+tevlnyuMfXDA0GOMC5PkMkj/bHI+B7T6Ix/MMduJ+A4IRUN5o7XKor4FjMciC
62x5tuZ/qhttwf2LDwpwmY5Kces5BT+Rq/i9ks+iy0NRyOF5TYXBedBsE81bvkQU
VXpUyVG2D83wEyHjWLS2c9sxhwjjXd4LMkfWKT6dOZ5weZezm4/bdKzQCRqTFUET
8E01UYY0GeHFTPnB9AoRTmInIe9VR1gEhvTIvATtb+KA31ioJQ/73fpLmQSAGQmn
bRozQ8ZGlD2jHpT1FVhRrA4bU0J0fFqZs4GESX7oF7f7g5w68T4K81p6kHWumD8i
TajubK2J34EYlruCC7c3SDq5Yi6fY1dK9ZjRYXGPoyP/Ie0YiW/gQkGbRS/BfYs8
f+dUdMCOsP6SWV+RRvcy7VIwUgf4XZGfQJ+xS3FRm7byjDRNJK2AabKk9GQ/LKUT
jqDOswghEV14vHcs+1MRo9deBM2dGL1ZJTQSYWmXuzNv6Krg2K5Rd1w6oB26KcEo
SjVUhzpy0ElVY6IRvsYsIU+GCb4XN8vou770eOGD/DXyK3nhtPnWRvdcH9AUXZCS
ZWW7rqZnShy4ckR0m7T78Eg7mYk0kIQSPNIZwHAwgTEOcF330Ns2HpHt5B/rGu1g
+LP13zwCPs0tfbdFvn3wC2DOVYAuGx5us/7KI/L7qagRGWDUQfiCqgWjd9tjTyBn
WEVN/DA9nwm09V+JcCMcuRlXqVOY4nLxOGkd5xAx8Ti4G5jR/kDYg/E+9AMYv8kh
YjgMZQ4U9buZ0YSXDBW16oRcuRByNL7zPQvPxQL6n59OuUBvmsGefW2Dp/LLO845
a/YtAx53JviN5mPXNOALTY6RZyW5Xo7xVE6kPs6NZo20so1lc0qLKtsLjF4IiAd5
oXOGFxLcCSutNPWZCZAOc0E3oQLXe+ML7EQFQrimQ8z8yK6RNxOMfYiiYzdgzdBC
uklT1ts5WIhr8yPwsIL0XRXvThcey4qcf8r+NT9JWDz24x+ju93Xl4DfAb31aKiG
WnlPQ+xca/OpEQkWnYa6RF45a07qstrY6NtnN/B+W0nTuGI9jC3Qwht7wR7KCvMg
vBmeRcPx6gmCl15nxBhlOfuAC6Ke9RC5ppUAaET/2d+vJayBtN1wh8BjM97ReVXf
+159p+IV30eTIp97TF0tHVKnVpMY3PE8w9K6pUHV0opn26kV69gj/uyvzMx9E6H6
YwNmXaMh7T1TUSPRbECXZx3MpZiT+1Uri24fZmQNmaT41HJEQVIP61qDycvGZ+bF
bWF0F6YAPxY4uIjARMR7h8ff/Zxd9rRZYEULDLSxpBa0MKZ8U611sPkbW4xYcVVG
ZnR2MkvcKrRlArdPgBoh3SqAJAe7aTx3/YHLiBdrKjl3cUu6NbOb5icp99BEYycl
ScEIy5XgvSqAGZbNzk4X6W2BrGQQrqdNVfxXHK80ooHTodPoq7uJqOZ+qBlCHtcw
8NHg5YFKHcq+gziEmyZTjBo65aZxbhRvirUfddAPkvwpKPr4yiLYkRHCg4zirjLG
OgXnEdPNLn0sIaUeS+FtOhuJ5aBXJM2mguGbPboNGGtOiqLqVpjvIlzRANodf1w4
2FNye1iE/oAcLaUx0Zbtl6O2I5XJ9eTT2cM6kIOsnLRExYOmcVApaOm+Yhv2eeRT
NXF6Vicc6gTrmJCBR/V9jCGMq4uUM2LKTRFKybEIVso6RU4SeRzhhzRRK9DymEcV
2Gfy4kquowuT+igN45J4Dq8jcbsuHVyp+MQ3dCmneA2RgRYIY/9D8iG3bzG1pB7z
Kup/H5JA2KS9cEehQ/Ev2hWUd6LppQ6i0SWt+sn7BB77nW2jasUhW1n0Q+LeVyJu
hgjkG5vfoKmvQMlcZ84b91yqmxm1E2jf+RkWg+IMz8al9WHKXA5hhygkt+CnZGhM
Ce1V97UO4QOxBzyFh8a+3D/o1raq/33d+gQ9ijsotoNTR9hXnThcilvsLe2mEtw4
CDplW3S/aOEuYrHgBuLlCxV/VDJQMwcYWD+FMfjMA7aaQPy0DWB7FdOgXRIa5NJI
VGOj5ODC1D1Eyv9zNa0cHhk/n3XZpaxfnB46QtHGK8qkJ+j2eHVGfDRoZk+eLpC5
kOzES4RmS4QXjAHV0P95/3Ui0V71N2Tj1QnE/Vjh5BQj6QWDmc218QjXKk2rFzkY
8CC5HHLIhSxD3Iy8aGObgQhuwOYto4aVly5ZkO/YHz2D70cFy5ePlPHFzo6DvQe0
SzGMpGhKj1ZmdxBH2aC8cUyLJcmIwn98NC1/RXHVqydgj9B9hPhstQa/hijOOyMn
iBgGXKqUks2GnU/TWO7+/E4oxGygoBeF2uRzuk655XfJNkcrByz6E6AxpOSfd3Rp
k7z5HMHVXWCTumDVNPDkJok4SJ+BbOvgyN2zw/G19FcsIRRWVTBUDV3ZTaaQOiaW
VcUcKX/svDa6QkYfwQyW93BMQmWrYB/X3JKBiry48wjagAswj64Q1WzSzWlCBqVx
SD7N7tIMuwWoDY43ccPRNF+KHioHkLDMan27a2MvpxHZY6L65kiQcPBmG2x0p8hp
MCgdgJdcA93ZE75k39YQrB9dLnd3WD3c52ua9Yf3ZwIYYEgKNemYJuLo2eoc6Uer
yyJ+EEs+iY4gaykSVHkMF+q+Q/U3yXQ6FhWA1wDX94E8zfuLHaja+2YMkoxEI20O
V1qwU1cJ2LI3g0DNw9FXLiME0ycyCXbmxBckP1UtSJGOUgTssFfkX8uR4ZHiQoU1
TkrQP6fEbtI927yoB4C8l67wntJq3lUoNxYVia6724nWYN2/V4yI+wMACSgsHf0D
v30RBbPDJjDG2wuagOLAcXVNY5wHLyvYOIVkoTi/hj6rDZr+vcpDs2yInQkmO8Ey
3QOCTSR0R22JAW44lNaPvlf2lhsxXlVARWMsLJQroNPy70YKHuxhFDJopqGEqbIT
fRwp3CoFOdmvZXGV5Kemjj3YLTm95RnReYoTFm5U9B0TEOYUBpPAYGW3CH7hr87E
isQ2gS7dWTR+tWbfcZhNAS+M4yYujP7x2lJIdf9QHUzSiJ4pwRV8+d4TCMvtJBDP
/7mcvzcMhWYPM13UW8sjY8jwR9ZbVNFhhNgsqcT9wOAZ+NErWOQ6ksU0A8iW2BiO
OpSlMI84Lv/6l87Ygw+BSukQXzMfpag5WP9WfGHV8qHYpu2gfejfgPNd9RvadFs+
H6BfFHZzV3h7NrQDzDWGd9n032kc8KaxMMymS3x7zB6j3qL3Khrh8583AqWuC0FO
7TXM0YblVptZ75xFxIk7Ui/+EwIUO+7p303I9FGXJXuYoFnayBqrD+NXiWfP2Q9p
r+c6m9v1/OqbISz90IFNsbr+SiaqOdc5Z4aBCWQIFoGGPbtZx0Fky/I3WJTFNDhN
NEhVGt8QWmaSagsWPc9kv6MxQcpqBdvPoiUmwncQHVNuaQmyAfi16RUeueWA6K8z
hh6rrbBF/ayT3C+li2bLDI/bIy/mO2tIpLZWaPvojTMV22mI/r4bbHCA2zQBgxOj
5DBGFFgBblfkt2cYIMkL8C0HZv/2aK7AzTMxVqoDpiYyHCCrCY3/96Ld1BZWaij4
bdZ6QuoQ9feOHoxzWOhr53z46LSDJFhYWgis2iyisWdr4oZ1ezo2Sc6ailrKK7Vk
/C96rtcfxDA9qIhCkyDMSgOUuSynFrykg1Gec254nlBHoXknA0oi2tTxpbsDw6k3
aHdM5FR0vlCkJEFXbi6ppoHuaM6niXTt3lqdhEEUHsDSapwVP9fu26+FSIM2Ubrk
NSwzaXhy6OIkAfbmMyDWf08xeAmAK4VuvjemXPfTXsQO3IhnC/VxKA6LULZdQtj3
yVFb2u0ZlDfwv+Ir1sFa4+Nc72mp6Jj9Io9WbflHmuM17t4H2RakiUVqTF3Dzr4v
6nDQWKLMo+uXGvx7EGcE9whZVfx4fdAlc3YFfLPfkhWZ1+Lo29pYx/vDGzSSQ3eQ
FN1hucpIc6bgVRDhpNN2YzdGitGmULjD/ZjzRDqbvXb0vFgHPPqLdrpZLBqeW/eS
R+cEB3cURKrC5R/kPMIqPvevnMUcx/eC+Z9QNz/LYWhzbk1ZMhL4V5eBMZdtS+qP
B/4Vlf1V285gLTMDEmgiOxZnEqaSSsUxybwi33XntM9/6Uvn9NN5y81x+SNXae3s
PevECJgGRgvXKIDUtru9960yj1rdxXPrBHUd8s4NhF6kjXPANJpj5CqjFsTAglcH
/haw8ho/adfMU5aTtbFgCnYSytTjHEw7DQutijlDfQQgV8K1iV7JnQrlgVEHDgX1
N4FH7feXOgkZR0eQFuzWlBlRYNQYM4xbA0738189j74dLWpwPdYWrGgGGNAszIyE
FaCtw/ddDLCrtKZ5lYiMDNGQH1FkC/lor2DcBN2FfaIroOtFWfdFPAk/YJa5SiWr
AtWuO6DSv08Pt0+9Z3kEFLKHTDxxD1C2F9uSU2GugxP839vRSBPEqhkct5eFnTk1
L/g4jyF21rSGTgRrTHX6ZXq6mkVm+A0IFc3ehLGVLrqkxPi0DLL659VRCYVJsyK6
Od1Bri2SUfLhmU+w7YyWpSIP3geXaJBMjBVUXQPlAVXe7X8eFaRDZcZ91A8fM7R2
07V8J1kxr9sVzH21YJw02vYhsQjPr4HyRdMLrqUsU8WGcoMXuEgNgjVEhNQ7E6uK
VV3EiMUpyW1+dahRg0o3X5kztVa/1Yga+pCP+tl5/zuGrg89wVPTEONvPB3x/1Oc
wx7fKBgpfLSgQMqFgP7TqWHmjq/Hq+xUwChHOI3g3qX/E4GRVcZmD2S8rlkBaB0g
xx2A/a/hh4TJ3W3MMqhoc+4Y4d3xYf8AfC0KCWqvNZQLYEkCuntdsdSyrLi6m/N1
cJC7/TOtfo3e7z5vFn/6OiXFMItV1UJKoGQsmlfO7AEgXLEGwluuOTwo8r+DIYrj
TjKytZIaf9tGo01z9ZSP9o8vgSeHOk3pwGh6GobgEJwrRFXdvnh2odvONPLUkQI+
PHXdXvQEA5LY82AKFHuYdb/lBVCJT74vSoi7XVVSL7IS3VbVSygPB/BXpOD6A3R1
HarYLe5OYSKZXwdYXMQH87GVRiFdLLUDSe2uTJmkcK+rc6zjziemu4DcTofPqnlM
oBBS0osoGbofEq+Ss+tPGVxqQB+pTXeEFq2jGTD3KTra+yrn+tnBa8EsiaVh7I+x
YCr8i8dXYfKgtM3zI1MBFvmXg1bm+JCOvN1RuY/YrNBMv/KWiU1UhkaghyhXfAR4
obgBOwyMpoXDDWAwGUPukh0n3jxZaqkK/M5j+K1gL5FgGxBF2BJRCksyYlnHcC4C
WpIODjQ9X/MWPCCdQL2GCozhpmQRp6BKZoTt5rpf7M4A5bIorqsrpYkS06AjAO+E
hAv52IH/YPluDN7VOmb03rwyjQBOiAzrO/5LEz1EWwOdkLH4eCTo5nNe/9+gPozF
C8wZpjEVI37Bx3GV2BVDpJt1Ckt+HW82+8aEC/PD+QttESqegPdtPHfJA0x2yz8b
Q+pazW3cZPH9MKkOPsbXo4EFCA6HCZZp92H08vO+ivQ+Ik4naEAo/JhGrdjT+ySv
mEngMoMWJftRjK6w0SFT/klvFiA35zJEC0AfSpF82wYO/7MYo0g5Oc3ljk7lb9SL
COxCxJGi6JTEf8nTURbeBPKqsORvuVjNqQ/dHZ3icvXVcj7T3ojXFwYQmobU++45
bbuLkNpXKloxr+f5ch3DxDO5HqjicUj5pMn4SspLzOfX35hQ1/gH0wPlR3+kzp83
YAQJR6O0YwdCggkTOqcc7uyKF0sA9HJnUWeuqQ4A0flz9dZpaS8XzZGWo6A70Svx
vuBldZhMcb3u035e2CXfmjTm3mOrJSp+9T5SNSTBYxme0KbIPdzXHxFm3lBRqg2F
s3eKrsDBsj66Q5poKSLUnTsITmLggTuSvXApTNsPhIJxXo7OMJMLbUD9Sbw0Fpzf
5U13RtP5sm/iQkOs6AOg559hSc/DE1VIomXXJFz5iqQSPFxi3d8U1+CQ9GhRCWxJ
sDpeX0fTLV2sxTp7Aho0asNu6UK6HfVOlebyY1Vcr3NQ4w2+sdrqpxaV48Pcd5kV
4NIiPf2IvuANcBCjb/iNPxZGqVr5uMytIjwwb2WSbupuxrO1LnvNK2d5whhwXFkv
xZ3pOXkq/0WtOeNdOri+XQJs+o9kvceSHyw7O9JAuPpmlRp/j0Z4//1B6N7pl0a/
8M5FBAlzKwicjy2Fj6f2bi0BCwbsPIzNIK/1ekzRnwYpbUZ8MDxSSi2AQKK+k/Tf
wog/7ILTOwGNlwvcffp/HDefsUWUNXPXjezP9GkEisr4NSuy+D3jL66QcrKrtAql
POGYI4NGAsfVulGkzUrGTQASwd+UzvydVAy+3QvWs0oFdi9ZMp1jfunPAKdfs2DT
yezVGiqL/oM/R6On4IhNUagSL6g2dLKFO41tFsfWHy3SqBr4SF1gqs35yUI7YNF0
h6HFZ+QGXhinCXY97ghPovFy2JR6frSyGxcy3qUYF+ptKpR/oQspGsUKma7Pfnj5
pBmSf1+ezPu3owX0PFaoZZzBElr2Yi7LznVJINtVsrmghIX+fnaEOxED0/vcCY2I
0h0LMYfSwE3LN1DdNM/gtiDsNaU9gbhX7x5TPqckdJGqUtl76CyZxl553DwzDJyo
YFE/eAgsnbS9mSUd9wvAXLqeF08DOJc7bbKt05HDIVg8yZ0n+iC6uRN89J5aDGmc
XdAhMrDxPnhy3tiIeAZ0g0bMhljhcvC4bE0eXTeGn8/33DLdgP3jXi6+27P0ds0n
/BzOvOqdAexxeBWZ7QlBZegoEMHaTg86fwg/JHbgvdtYo4JASIBxZbS7kW81reQB
hcesmaiP18Tga6PdCIY1mYHiqbGjmKCx2Roe1svKkb2v+2OEw17kin03hTC4Co/F
LPI0S2dsksGHh8Kh6jAwhZ9HAi3QLhuB+YTTyIQIhSzc21JYu1p3WWsSjX9o5nl8
z8OAKCmhL2ktIOmScjbGpoXJQnK6lTGRS9wqkz05Ru0qjEazw/ZsvyzPadmbjZ8K
5nyxt6QoyvHSbwvaeGo+TgJUHJWa3TWLOQdZskFLh057zRzqqLaH1iBd7qQAdTbr
jr985gNIo10+IJXUDWjuMouALy1cRImO6oipABU0yE56nHGXKfAoSAzwfaH7Fsed
CV5guXdyN2pFTkT1bzaXSRY7Q6NHLWGQmocpnk7EZWY8NTOtIFcKOvy2CN0AUQZ1
Hlno9cArc3Zlbh6/qf+nP19C9aFz5Pemo1XbJfAN1Gzjg7oKSGJeKXxZC378e18z
WBNI5CynoFeRB1lJk/zWT9Q7/gwKqrkpOkG8O4OdrgCW3xghb/BQKP5TIcUx6c9b
SKPDX5n6mmYXWXnMntj3XqfLoFx0oO3kYxKKlmWx9tj6+3xuPsOoysxrCImhKoQ4
cneqcM+48FYVA5zVjIImqPt41i98EZ71fE+0cygsM4jcXOEM9W5aoN/9O971AQ5W
RQOHCsJArXtuYLOADVY5L93LA7Rh0wVDfN+pX6hhQXSYy3Q05x1XeY+gqET1QHwV
qxxBwRQF74iHiiXMyi+ogVbuOnAUPO8+q21rIXwYmp8Ro98maC6UkAHfnazVLgoC
44HGUPcI7WfHYOoSXRs/kRvrGfVUgpWptsN/vMYbmv8tXsshmFIpuHXHaoB31Z61
WNnAWI6EwSbyGNJ9p8+3OramnumQEpnGm4kgyH1/U9i0RDyoFXqUDx6qoURTE9H+
F2OdmEv+FAWoMd2kPPTSjAtvZEOqLEin7wZpV2IvH4G6aItLQ83UmL3zSJv/BHSy
R9jAbzDqldP66AUHoalhYLkt8G13+XYwTgqhY68GCk/tZb3ELc1V+KcSXnHMmDij
NFYV9g979FDML0Zh1oEmDkJXzLCJBoHDUcu5UAY7Oo/m0iOap1Ou9X8hYUi80b/c
D/2O8S1ngwywtewanrDc7hRXJY0CaCwRB2DfSg6jmu/7sJngIKQBiGj3KOq7si8R
g+1zeqYA0Q0POfNUz9+Yz9nJcbXpfGpFKr1XcQUPDOJapB2YA76sivYMVpPpi7xG
qZATmQKX5olVv1Lw7efOjI5hatmrlr9rXvW1TH1bWZe9J7zIvjPx8e2gkH+9xU6Q
PiSKwoXPg0/fyU2NlqSy1Bq5oNKB+iT7QIOk+1oBUsMc0wQIfwIL4QSf+mbX5W1K
CnenBdwAkWYP8qB2H3hnf2Q/Tq9Eh0oG98UYFIPn6/wS9OsLF0yhodo0+pjTSqZJ
/yd/AhwuJ2Vb1u3930/CJWKK0Bezjjo6aO61cFdwXB0HrxHKq3laOXO17jbN0MLu
In0LnRzAmSrBNJVY11jWH7fYnn7Y2sMKciXd3YWu4xVZiDhTxWoQd6ZXT85Aw3cA
qfy8rf71B9lXVbpvuV6duhR7u56M9jlokzNj81HfAG0toqkt+vrQSLRwlEf4bntR
9IEcOHf4j6XVRNe5c67IOlwpEkX6U7DOk4f51ZjORv3kff5pwHmqidjhvE308qqa
LkzEVsw20FfYR0SBZL+W/amZniqx59BT8iZ7umchuOXdsRt9Hp0gUqn4dxPWZtFP
CWHJqp7unZyVGLMKPWfoBhtPsU19ag1L4zQD9tmxL/1cNxmKz5CMUmfbVs8gwmk2
V3pwkgs//nAs5t48gMZDLRRFfTBeUGYdPu1yy9DjAqu9g/428XGBtewva68Wcyvy
tasQv3Pv2g/EYX4XrLq6V1qMGL9G1pcOBYu3bUyyVAfv9/A74EgSXeC1mkEdqvFj
D8B2S/kaSINMB8h/LVpTE7sHATrHO4w/P8gdSv5oH8Mw/JFSfy2Z9GdpDoUL1/lB
t1KcTWEwC8y1nw12nTsx2kq0cg7uckqJQd4HNi6LGoFw6HT2TH0ppZdzL+E9G6+3
41JBJM1mc4IPjp033SEUMR8my8vOqozXDAcWpt/qufGc+QFS9CvxNshlGr8PlRFZ
/KGjnblsvtGMNbh5oOZ1UkLXRktRgcgerxlOuoedl0EfGanQpWuAyjxYg96S/jdS
oO2/x33+nsypSoUKkA4TcMcCEb3zznGKD7+9DZ/39C/K/9a5m7jgZIT6ZZOupRJd
LAX/z/K1CJ/C0o1tviRCQiFkrob4tlcpCf/l8E3yfByDE2d3B7k8n+xhx3QG32pj
d7hjLmpfolBkJ9TdNu4ndt/F851PB/UB++80TtmicjSUGWpaY7rv+SFBk3RbRG2v
cRi5mZJAKsG/9Tqqyy3aV/IOrTaDBWXnOs0fr4OAdIyYwp0/bNNCYERI4f6u48Pz
CGRu7iin4nuu6Rfzfz4w+3cXAaGnx/figS4mCtd722PJOFKOv33lBr0/NWIngOd1
HspCNRFFFKC5uhOW4MyVQt+O0P1xwMUIYqKxJLKZyVluM66boa9Z6NyaJ6u4fUuN
uTBeGvu2oU79z9afuXZDKic4ecyIzeLi6WyiYwng/vf7v72jfl3IVDSNMsv7rO/I
CHN3YquhyPSzPgfgNCwY2DCKWWyDQirCH9fQtoys1bnm7isv16aCAHvi9B6jpgI+
6UkuyjxGELrgnVk+01zmD1d4a3Ifgt2ReJPDu9vEpYIsmMOJuIWLW1OGso+c50pd
o8Cv3TQdazuhDTjL23tRMgiDLdjWgPpsjx4kSw6aGPGf0kzzuMubpHc+KL+Uceop
BJQlbNY/uXKN8TfnCN0fw7f+J8gQT0u77pcKVnz9HokwyJCOF7fzDgQNPrgmm4zL
oG8NyJzg+LbWsa8bhDqEph6SNYWz6jd+EPIxdIs5Yie6C3ATy7oRR/9yQd79duvh
934rKQ0cTHXurWPTVFi4RJF8v2C8KaHtoZpxaQv6afobD2B7EagOXn6ERl86RAR2
jJewtbPKX8rCxMhm1CYfk1MFS6r7QvA3pQXqjJJrnkWUUb2+mFOJr4Vfjj77OE2h
EvY49a2i2YDO68sWNtWRa2+T0memquSX8mfznjWmdU3O8Dzj60OFN7We9pZfnLnZ
t2A7PT6LEF9hoBX1Fg8szMLQWB2qqYUPo9eIjn6s0kQMa8x/uMUHOGfpGHjGGMoe
22iC5VGS38MwwpBiPe8pDpdiULk+rjxpKXSkt2FN5F4YejoWFdf8X7ksK6hiSW6u
FAd8/++RD+X+Ev6hBJ/WH3W5N8wa7pPq/QtcKsbSVjXRtNh5aPyPjpTPhBo0QBem
+Y/qtkV79J1C48y+utvZXnqQznFA8FQUZGpGtnPY7wDaZ8gl2sNjLUgwomXWJ5v5
O6tMUlxaKqZIt9yUg061TF6ngzHbU9YW93sKRd5E4xQDsuTZ8KOWqTNoM40A2PM1
/rc5zy/fQoLTms+W0AM3T5I5/ssCCX6E+n/F5wd6pAJcwBQpAB+5c5jR/qVokTjv
HeYEelWQjGJf9G8HhfoG44mj60rcsjHZVQAwZpe2sXz0hUO0yCjevfdxls3aeiIb
BBlkIrPZ2wuPqkG/87/dDSUmQzXmFrnMxXjvfz73EDjcVXAmae19JMGMeJ5rBai6
BGklrcXtktT4A4Z4FkRiHwmrQXtebMiTCq7/tNFPdkP7FFImhl6B3lF+Jvout7Vc
bkuNmnn/FuJp/ksN2p+0eOgN53pVVFibzzVw/Vy+rm2SNws8MHII52xkepKDqtRU
AX54gjcTYvo9DrsBMQG+AKEuy7mgUjVYgw82KvOGV84Py1o/ozCweSlTpkQ2Z7rr
bTF/98hIbbi3VMY86LWw3wjQ3IsDOwBjpSnEFZom4pHDHoweXFGVH7lj+jLtKTc7
O9ty+CHlOBpXbV2RJZqjZZoEBFVUqRihQeRGja+9K6RTkm1+KvqOJLHhopPGrXL0
ySEjIiW5k6LJgGZo3z4CB1I9gA35HUXlRIHUOa4Q7aX/fkWrUt7h9/rENOfkdAmL
g0e9oN8DF8X4IwPrAv7t5JznQqcilq3FEvwTtyllnXwI+nSqGePUNv8lBRKYvh0I
D5Y4zEvUhJXavrM3qSuGOFzwzD8vx2HIrS4W90ZlblGZbdn4DFoa9ik73igDgcJl
sfrKjY10BrI5VF+EvXJmkJsm4vreVX+RCDsPFapS6BV6WOA2tdQSaLS3+BTd6iq3
3hKPZVk+FHKxi0pyopI33Ykmzyz4cNcPe7QNvhlHX9kw91cEHAMGCpSHFByADva4
GZ/hmkGquykgPkBakme5AfL32zc2W2TxDdq60fDK0O7syqa6qTZVZIsfMjsKimEG
8bk91kvMgpVGLkr+/niNNDclwYjvAtsJ5Z1CymW5p/dEoktMX2EGWZPnYBuqXrDE
Gw6NztLA0bZqzOlZxC10fMUS9ZJ4/nbSoG+B+jVJFJD761rg1my5/LVayx2jAPBx
aQTNShQ0lJd2QlXrn2AP4H5itFC3WARZdawMVYC+XidS7kW1dyu6VEXKPH5ne5aC
Oeti18T9ZyO6BFbEnuFChbh3vJHjBhRycq3ay18qOlXZpmc/fYeWR1Ff7U1O8Bfl
EdUBeoq3tMsOwFiEHsciIkjMTysPV/DiBQPD/lExlKwNjqYYGJo2RMLoJfUeIuKi
48QVFco25yeRAk1aksbSeKtwPFDN3HXgxzqmTPodXKKn8FMwaOc8xD5xa7k6d0kv
VQw92jkhVvG/X9vS/9lsSbkGTK9agqk+Dr6xW+40ukiAakfuC1SC3OzS9dBCKLU8
n9K2SSgAdl0Hj6DZW4AXcSB2B2RHM23ufxdIywW344BqQooNRx0hmvwA1mTmSJxi
fcNSCrNYY3MDWzkwIGBRGC787aw/RpUrwwk5Xu5U2vnVDBHuqSA9QBGb85DGRt/m
r29zltOZUYvh3PTwC/DGfN/KZ9HA0SzEeyUbb4taknYt+cAtXaCmmUaHzYAnC5hN
31uIAyoWAhF0sn1LLz/u78UsaftGvOfOECbTwR2fPJ5fRUtLrBXSiqDeqUTHTPK7
RfSq7RaJ4qd7mVZRi8LtR4E7hnDXnSSXw9Neyg8u2cflAfuYRFGJbO9c9K6RMYPb
KF6ULyvhEVkL7dbn0Ky7RNF1SbAdaA/qqSRKlR9DtTbSq5cryK9DnE6GePc8xTHr
Tk1B3gJbiEiVsItGhS4V7sPOPzBkqXaWpZBiG+qPV2Be+ZBQ/eRyfBNFNsDMMBsj
R2wnvU2D7VKcTsUg/RpfhcMg57TCwNTI8fVimDIPFMMIfTLrPpcyMEE9uyE3Eb1+
EG/wQnIIoyGGGBerjdRcui+d8+P1mS22JmKGV8jjkYB39Gv37aNMZVbT+12hOECk
qB4yKgCt8w5dmaJUrc+x2RT+vdn1ZvgSrQMBP9Cl/AXEgeCNrbgC2QTUwiG9Jweq
ZVf2d9MZ1Ea/DK3pok25aSxQ5JsMqaXd4bLNVcM3dIAahFpwZORbhcGIySkhMVUh
RLLTn0N+WH+JXeiz1CoW+G4Y/zGgwfjtim4QCdupmhhMh01DfOpj/nPE+eU0HAGu
y2UxyPWlDAoQ24fS6Snb2W2lZwWqzU9YezqXKJB9cz47pH/qUhpTGA07a+b2kWZq
uwFMEo6xOQktg88ZETnWoSv+XOj+Z30K7FHXKsrVn6ixsRRld/9TSq8BuKa0rgM6
bqg+OIvE9rz9v1Rf9vFSUOK9HWp5x/Nb3DimLQtL9IO3C/t9vrKI3BKSKNjNr/3c
ADAR4+BXj+wK6RS0EmWB1Y/smXASJB2DsLmvOoudswItvxmN6Yn2luMGF64jcHin
JeBqFZ6OwNUrLTRM1t/sqEA+FBcDoSHVDNVPmdnC2/WeD7X34puIBQzeO7mmYRDB
5Kw08a9MsWpHUDJE46x48ihYiGjf+N3DtVuu5fcG+2JRLNuToiui9hJSthx9QIaw
tphqM001f3b6YFIb6YkJgGsbXzAEbi9M0kHYKTqe/kOBrCQPm7iC5X7r9iOyv1Wk
BA00oQNI3//wy+SKIF1SRB8Wo6KvF/k8Hjo1rUJihqvKck5whr2Z8bZYX4jlgXQZ
LP+yfSNC2Be8AJtiPb5ecHZVwS9ivfzMBC1yxz65WyEpzwx1iAxCoZKf2r5Tef9k
H92gKp7iQtOuIoqRezXDBlI4dNlJ5YQ3dGXfFfm17EaU23ahZjwSFMn3dsaLuZPK
07vVlanvu5xjygMtAvo3wIHS3goK4Adv/IlcR9g745xlYWbsNkn33C+Sf/D5o701
ssxiXy/n0acMa1n71srSWKTFKz3NC3V+/w0E1yYv4/e0TSrK4yKCYAQHjX67LWSF
g7vpj0jLpUkbYUEacgtOO+gTMOPNJ89WGy+JzGHaPUm5K4X4FrpE8ltVb1E4yMak
WKx+AO4s0LNmBrGY8d3QMYgOaopv27VCP9p1l4MIgDDLw6m2Wm8j/cyVr1aRPIzJ
3Ek07l6cmImUZv2ccgbWJ9Pmd3PoXEuaYmMQ5Yo+Lp+ro5R41VyTZ2SIigdwoiNr
4g/HXKoA84fiZl71bGE+d8yYCxhp7r7NXgeDKAXGAAcFAZsrBrU+398dcz2qYkwy
MQ+kue763KSBFpuXkHGhliURRyI0lhgT+jZim4oZRPZ9aoJb+ap4Eo+fSYmjBNs6
xZEa5L3u/KP8eI/gDwfvjvslJnc9IfUrKhd666KjIuZAn+Uq0MiNhjT7VsgrY2Df
OWRRHCci0VKekc3mLxDcg8b4IlNopCtKUU+6r5sfU1Lq482AIV0xTWBIH6k1ZDYz
BUaGRwKRhvDfRRwDCKw5f8ya8nndEaW6mSe/SXU3SALktXRYc16zreTxnFdgmwPL
3tt9/W9jZf9fxwMxCaPAB+vUY/wUpUrpyyjpkyLmYEm4Dy+Uw4AmYqUjcm863jpc
PczeoNeTKrpKc9cjThpC2KOHe9TxrgzVGMQrg875QUyV7qSq42wpJHfdi+ZCocb5
BNcxws3/YSgjSWiOZ8TQ3/t7m3Sab+oRbsr2xX713GZDMj2Q08A4Tqsq2FxhmsBQ
3WE5cntCEsvIOglQsRQZKJm07eSdxNLyt7TRywH6JLMdRTx7v1+gSva5YcA/S0z9
gH3k09L6Y1RbnX6r0LrWd2KEGkqHTSvaVNHiQQ6ZPwiAWJotGUVKtUgeFpB7KPfA
pYtOK24mZ9zAEpq42UEageCmimPDu2YP90MrfUK86K55aXWi5tybFAJX4FBsiutp
eUcorYbig4mw2FS836uNJ6CHygTtZbenn8oK3b+j79V3m3CU7OrnsfHEp/edqH5T
3ExUG4hb6tpc2qUT0Df8v2eyTGMdJaAbgqrihGz8ENUQVm7IEOe+Ns3S5bR1sxF3
YCgaNuoIRI+h/Z39MJvHn42ntGKJ5mNVYwOccuwdYFUyaRGuilOKpngzMalhrZ+5
H7ZeVSzN8XzF3a/O8LShRlv73D0Z5iVRzfFw0Bnt67AbPL3TyCPTaqYEPjptRgje
43ZVMu1xofw+8Eisf2kpBWjfxDva6wzxG9Rnwrg/K5HOgUtIkccQqUpQFpgHlSV6
bSgUh0Avzh47cr1KKy1rO0jQobwfwD78/5P0/LEEeJiEJOOhQPimh3xtCQGRi1W7
ET42xDkm4/PfqOqjJKumOKx+NY/yfLcjwFREbRA4Pnd7E3oho4eELvxhV9hovc1f
98tFeT08dYcBxw5euH01jEriuBotiVcSoQZP8JjGorj3Bc0Pz+Mhv+0vrDlFX6LV
Cf+sNCF7vKs+LyqnbcDnU5WKY1yPBJJThDROje7DRm8uHfvDzKlyL0foU+jSnv/s
fleX0Wa9eWML5m0uo7BelhINBhxVH0W+iU+BaOiAgGHtIMI/kWmIWu4c2CZHh1A2
OxttW/a3si0EUz3FBdoTOAgQfx1v+Wd/Ra+Jr4OtiYItbsqDTayRhZJyFysWRjmJ
J8UiLCVNJMMs0JzI5hWHxcWK42v+rfIA9z19e6ErjHeVq9PLdrziaS24HQDc7hil
Cf7jEJ1wWp8/XhbyhfCgBdOJaSIRrAEMCqRdgyORA1aHH77tiW1p1lX8kRdoCbME
1k0OeSpBmUYYYxaR+djOcLy6u4pPOFWyo2x/fSQOZKbwvtVo/rWY4YZ2ERcTOjeA
tw/yk+M9Ieep9Io47vRbECAYsP4deA66hwCSnZQ40gdQ+/s2al9iu/Y6iMJENz7q
i+x0um8k3TgLjcL/3hF7r0+Lz+1EP9DEfP2hC0GU4q/ZYJ/lp37UeH0p6161rBug
Op/pibMUTW2tcXRSQwC3sVKWHwNdwDxE01ieUukKy22hJiB1MXXpl0pBP7dqsUdq
Zu5kqutqc73lbRkyoD0CyPBG/2rjqrQeVRG8FZIZjbfUl/G6vPZWLFi3VS567Q5P
KsMQBDX2nROztFYFWXukzmQxydz/7/T6tU5H+V6q6xLzBB5QSkOebUYOZtwoShLG
Af22crnaSDs6+sclN2NEkBLUrGXXdcl1otp89xxTemrR/UHALusQkOL+O/wEYoJ9
yoFh7qzznN2EVBS1oguNJJxfByMIFDI0xygLqHaOEdcAUhuexN9K0etf+l1DIGc9
aP/d+D4dcm8gbu0HA5dFYVesPDrDBc9TGP3EU1ZHp1RrHyppddfDqgxbUXw4MC8c
2cMXHnu7e0yJoAkHJwAkEWQpDAcFgG0ALRen1C/fc5GeRhUZmWp5e+6LVP8iLSvL
3w/6F1vTJ3fHbnijGBSZSsFB6T3UQw3iq1ddFOxR5oZcLF6jZ3rpnBnnlI6uTzQE
123V+jLyzcgnf+8QVsMGgigEUY4pDus2w69Am2lP3DQOzibQ7+oYZuEW3T3UMezV
8Tm57B3CshYch7blzW7WVf2fYj8X/XFwj09q8E6wNG9ZNyYbDD6tDmBc7liBkWy4
/fZnyRu1gJlDbXTfUS2eauJvNg51lH7LffVk2+0mYJXy3HjcZKNlnfWhUJzfIa6N
PA5fCg4Owpyu6y+Kf9wVUyJraY4A6pPQVvgX8pQ2l1kRM6eqsbdH0DFgUN4h+uyD
srYS5G0w0eVVfP7l7Yh5LJWVm0xSScuvCFkyqPQd8jWnxlhPYkszaISVWF6NU/w5
DBmS2MQ+58exD1DoBfg2ZVw9m+TVtfAN+LuLTelS3f6fqCg5P0Gapq/IdIGchpxY
+5ut8gNQc1W8AvYiM7SAKlMpvuUFr6g5Nv2Pg73FxQHflrOnj9NYDXnK0gQD8piY
rUyb7Qb1QGSZunofquU8rOipyZoJc7h5TE3LZI6FIXNB9xiZYszyCi0Oc2QExUJD
cLjY34Hmz4EeC5kDS4YJjlTNI08MFE+I1FBP3OPVz/cE7lemKmHFeGuc/ZDgvebW
HS09PXi0wfHsSaL9zsXzsG+OGJIL0Vlkb4gfCrr8MGWfdD9iMiXEnHzgysJvpiAT
XzbvUy97bfT8hOeB2Fx/b1S7jotXcvdh23Hv/NmH7+ntsaIX+sIk0IxayUVE3Qn7
4SknSKGv7Y/KDcVLwyj8txKGsr53gJ8X/gjS06qeZMCe+P79/FsrMdP4du4uCwxZ
GVPQW+iYECXa8tlGTUVo6OcHw+uFFV7PX9+MSGnZaAwAJEZ/kfaihdyh1rr42fUM
Z6BeCwpsK8OiyREhJO41ZauPiTUtTHPWJTJILfe8XPXhkapNM99UeaWNVeSpqlyk
gEtvDbX8nw8C6Gl5okcwDpgmWnSa4BJJlCgwpzp6xxuDU2AILSXCxcXieYjTkt4j
+EhMZGXs8QFeFyvY56B3At80HzL/joBKyA4pIJo2jRqWSnrQAdRaunU98eYbtiOH
sJnuR4x/Gr6NqhS0i2QJeqxYCQHALKllQQRRpWRQu11+rvLG4GjafrBEFKXhHLXN
m+grQSS2invWBfz/26Nqo6enbqOWGtAOcelCgGpvbsLO0pSPidh++NuiLpNJfGOj
2j8FKBvzghxQnb1/HipeqlDSs79urtWv+6pJ41eFW2gO4r7wK0JHHfkjdaEFyA9f
P9oFpWCtMuMstNYaRNwUa4eAzGDKXo1i7IjP6jrJXAg6NMqqIIoo8SlkdKol74qy
hEQQ4vPezinNkVOP58Rgnsi/IWbF87VKgcggMKcCufwdr3CJwRldotmgD4VFkZDa
RuC2fUQlTXivExxM6XK6SouJPjcwfz70yKKXpNEDs5hhOk7yIv919b52r4bAzkuj
9JYM3fSsbT9DGZJJY1+g31n+opSF8lx2F9HUc64ptP7t3O6ayEdStnBoz+lZ5jHo
Q6L67CBFSTuXYbNS0Jam+pVbn0fpt78ota++UywLU+WDqpS9eMeWTn27USmbMy1g
Y9PQYr0jtcvtTavEe/yTPYp3MxAWnuFSXGeLX0qPagaJHLw0CD3A1qTdq2XF4zC8
q+bAst1X6hoMTqf+F1+u3AQwPq0p4RIIeIQj5d/CNEaU+olpEYF3HWdoiv6GnK0C
bzWuaMudc8xKykEDSsgXO/2pk1qLiv7pmmJyDybOsTy0n1RKSeqHoBw+S60K2yjV
vkTEodF+V9N8Su6mQUqmPMl5dYBcO7TFjwjMB9JZyt8XbN2y80rUQ3u2J6Y4lAG0
nhhiQgOcFRWyee8I4pW1Y05UatMm3wFCvSvtYv4BF1QcDQnDIP1nLJERNTneyve7
RGTq0cveBABG5hfbPvi4FoLMxrGPM+YMqzwRZ9zVegXBY715Gl33nh8pjKb2oQaU
E/cUb0VY2gSDZ+pcZljSX+q+L/pnsj8BIOzTxS8itVPIyiusU7zfbC6D5Rbg4I1j
8YCJfFreGlZOdCgS0JfqOBOTGk6Fw9LfIXbNODK+YhNr49Voa0HWR/qAeg6NNVTN
rKVu4NUCINbcb2QwoGm1SPjRQMO8ZJzmSj+UGNHVl+CaX9QR4/tCdq2mMTMGKaZq
Tbl5YQCLOCXNiO4FqEj7qHCfzJwRVeyLApGfQFiZZDFvj2LfW7YqAov29OUSCuXr
v+ctmIz0DeRCT2gvmlkjO+pktyDpTl2YRGD4N8pv4pwlp8EuIRweSeNBYV2DKlV0
bKd73eIa4wM/6NtIfrY/pnKuKcPdl4whjhzbWl9NtmS0K++5rAlaNkvl++mAS3yb
/U6vW7ZLXbggcndwyGQeDFEn1pA13GABIZ8QLBtzl2eIPTW4Xju31Eqt7N9fFZ4t
me8TSjByUyJUcQi94fyPQQErrvykuzZviqFIn6tUOL94dXPbfTcCFUKPRfU9ppP8
y+Jevx9RH7EIR6Xk3q6ZbD02ZwYJdX3k8q5NhWx+WwK+KUHoWWPwnMyK7sQ4mwDx
4TRg8KLYVEWumR1s/ULTca2zZUcPYUsKh/nLfURSl4SBETdKVD7UqpTffzyYsdZ2
dWnYsvXPJkN4Kaf63PbciFIMnNUUwPZjWNF0EBOnhcBnPTAyyjFiVnlmltBt7yu/
J3MZRShs/nr7fnCPB5hOh7Oo9lVa2c8vA9fKGBtfT87ogqVORORF1uNrpd+zj/u6
dfjHHCrvORYJsCt8N4NLR3Qg7bMpBh04f1Mg2vTaj7jdd2s19uCDVjv/T0bPHRuq
cvCqJjcq4BX4JEwCshpK3/F2roEXJ8xgZKSSPqnLPkusgpCqnmp913AKKcHNDyQe
69x8emqQwMJO/0oLDEXvHiJITc6hfIL4UdAost2KSY+duDmeNDWe856dfpKzSgkJ
QiRQD1/Nx5ZKnU6CvASxrTktbzVfhp212uoC7diy3cKfKhv9rqlI4DGAmxCm5s6D
4MWRCOSnBqEl9Pne9k+vb23b7I8pOwDRKLlzhBso/X25mInYuCLMufoPGeAZfljP
O7Lioc9fCU08d/BW56YhVJVhst8YbxB82bpw9K28pL54l3HfI5Q8snTJ8wGD9Ip3
FlHrLqZbwd9fENxrg5PQa2jDFcKtp7mOA5bF27KH60mBwdDPAqit/9Ie2SB5QvYd
TD6azx0vS7i6koECgD12AtwlQRyaBh4yIgAEf7Iay3KVQJnfA3JxwpEbKivwagbn
qXSZvhOosPNCabzfhMneWJ3P4LuFGLjdbdaSY7LS9ByY7w7uA7bzgz/goo5HAevZ
Fs4YqVv1Gj0+F0ZmdYkU9WkcBbSwsSDBW3FC6N94zPJT77G2Y7WpK1dmx/KD9edS
unZLRvBiyly/a/CY1HlENMp6nYeWsc1dZpFtLXLYOyekAWkxaxg/QtGz9K0R/I2H
2FLD8kjec3ZiqcpC2pOLSQu28dzeK2/6U7fPK9xX4V/KlsDKW2ueAS4+foCPLDNO
CAqE+DSnLsI3Q/CK0b8KVrTcxa5fz4Ky0cYr74XuOWbAoxyuX6VwX0MKjuyg8MEZ
HiFEPsx/yQxVDGyrL26AVZG/aDstdCA32lPsu/Lxri8uWE9l9sj0qkz1d6b7jPtb
Xzwhrp+ujHE1cABeU8xJGET3keZKc4B/2cneeyjBpg9HfPjBkkWMDI2+/oXmHc1X
bVSM2fkWjLccgRkMckgC0lCAVgqkNhIuNVqyZ0xon999Uco4OwrEjaVePR9E1vGJ
yTZYH9G73cT52A9m112Egs1iLH4ZyWgVYr8DDz0IQs9Rk6qmuknbOis+v4C3R4Qo
DVYu0zhRv+iSOopBW+bnxxozgadhBsKRx3jkilmdylj2OV5FeNb0w26YWRFxMlvT
GmPY+Dko599cKXo89VLD2MGrAGvaUCDdBFaN+2LV3gPJLjGFCpApkll/U6gCPHHM
GmECSRWBLk7d+/vj6NlCV6BSS82A21bAD3nk7SK6gH4EiiNTSmNvof5jb0ZXL8L2
45KzI50d3plfGS9hyX1zKRMaB8QDWb+xQWI0/gpIdBI0FnoFOoWA7uwV/mARrJ+o
jWXtOtQAFJMO+n8WYy6J5pxNF+rPiIwU0ZRk16YgCryfBg26E4mx2RlCrHk8HPy3
lAFlyfxp5TRYYZ/sR4L5gsFuNHYk9gnXv3VU/pIuEFLNDeV1y/TnVrdQQi8Nou0Y
+ZcntpG6bGtNcFcvd0CeSsRzIWazZ68wTeiFT5fjCWBYoMgI/is5oWRS15aNxKd4
XMcGcDBs32Dw95YkMBCzYNcc0hxb18hKszTZGZ/GRuJKDG3gedldxLBkf4Qcqhfh
xK/ai/8ixe/lr/81qZ7spYbBWUsMsVqguJ2jruC3mFzCthO8478uhilWmnT+YEzf
QQQtDjTJ9iGNDPEzgMClVX3N7ZYFtb2pLY+pqD0zGh0tfw0hcUz/xe871tna1S6m
KYSnAimOK2u2GZchrfD4A0AJXWjmWgOvbpg2tCgqzPgH/0yy63I4Df3GBRHNzR4u
t1TONAtLiffrN/lxE3LOYebdh7/Qwy7y1gA5IUp0ltquJoQmn/xWNrN1xljTKMNS
+k7/8ohNKOy9HlEEAHpPpzfJZVD7ACHMa8pj9gPM1ZA1ld6D7jDKnG1w60fZKkaw
RP4QKDH+uKX8MqwhDASs+Rticyl9iRc/AhlNIAUYNBoCCbh4s2iK35hjoWqua8ZM
02lEDMWUFBLyx2aFKVh4hqidiHEMiGGRYZmiixvqthpGRyTucD71Wx9DUABoSCtU
s9tv1rafrbas1mg2k1H+tfQvlB3oIybbI8v/mq0RS5lIF3n/1/Y/y79oH57DECED
RxaowSplHLttNGlqHcobnplddnKGQAghvi4r1xU3IVGHP6ha8POZNTKKmV+1drHI
OorW+i6HZb5KIewqBmDkJZYaxXF3nO9pXLsrrs9WGSfczuBj2HGhT/UiFONipLTk
5LB78xBlNQZb77kt0dFut2ayPfEb/2pfb3fLMNpVh0kvAypEENeXfvglYpNGfKyH
vcCX19/0U6qa6270skrRHMk6nC5jtzNxQnoNQEqZPNj74P2czmP5d9GTeuHcudqu
8RoNAcr0dmYg1z+q2xJTLP4MsXzk9q+TfbLfmLGQRAFl//DQcuBsn9SGnrYzY4OT
VQnFk0BnSjIaILlCCxbmCQnIJ4dT5Y8LK/K2kP2Qvo7yyGz5aPwvZB+3jjT5Z59U
1XmO4b341mSiZr1E+kHJfEwxsf1/iHTt8q58iVXttkepmhrgi5kfOCX4NLhABMFe
Agt1z1O9My0zAmBoiHWRmGHjMnJTv+KxAEhOyLTVr5eZqYvRO++ysIlEyIL50ZD/
gedsGS/TjVns8nRkzhOmcn/+gYKyD60/oyp5vupmdWgD8R1W2rOC/hMH/wAn4rw0
83LNzDo0e8WcImvrqqHSZaPC0gpif5xRr+AiqmHnHIMrTE7+OapreORCspWz9nW/
PUOik0vBivyGJDmD9o/xIrbpo4nXalKW6pJz93MFC48l1oa8Oz4CHuWxjXWYG6hm
Ccnsb4t+Xhbip1sZJ6K1X/4uxJY9rwrdeLScBj15gr0SDSaBPcjmmfekFSr86zbl
QThrtR5WAHCq/Scyk/EbtqzbjW0rvl2ByDePNjFrrLQpd1hcZynDBU44LoW0J5P/
I4QLsykOojBWsD2ImBmTkWctzPwLe/IYb3Bc/4/1ZNER2CcHW+1BKXzsp8R6iiJf
F3nW7PGdQc7AowyhficQ70zMTEFmeE/HxX0SsKEo+4FeA6iBd5aEmgLEcn1NQqqv
CrJTg4Nup4GC3jYnvxJyDHi3Vno94aIiodVPPNhiX4Bv2pqT+015LXzIIjl3kmyU
eVc339f2kM4Xon5/v85tX2TIZ4Cj0UZIapJNQq7f1ZYVLdDvqPAhkqBFj0Y8jkSt
uXvLw8M0ciTQ9Eec7l4b7saHSYaER/63cTBUwgfBZPyfczScyvuX0vjU9wuyNaaC
DuuzTTrp/HpkSkxWalYPx8CeVRy6J0uvDrM7ARPBT5hqiT8Q5rDXwttcBBaDuf7H
stWUZZjMH+U4VatFTxHLlzzH7kALS1kgsm9Svi0qURfLvwjcsJ+Oe/YS2b/sl61s
m/xBO8Y6z1wNCm/ObEmmly6DfTT/n7FaJXfkEfPFl1I2iDKFWdctV+NCGFbwTAbv
ggzeXaERQ/lqOthPJ4Uya2S3SsEHkYI0oShur5qKY3B58RUxhiOLUZ3z3KnNPTuI
lILPqY5qQd9AW3JJnEf+vFjfi8XWWTrDw2SmMIWNNgL/7fQFsS54jdlh0+SKzmze
J5FXp8BTQ3I3p2IZ4Lerzb38hAvR/KrPo+kSVplQG67+je5f8uUC/4yQUuIdIP7w
bzIRfe69hsccNSP5LCYJW70ZxZ+fDu1gP41WF/b6GNUP9nufhS9E3HsIU6meUM+B
ZxquQnPLpRhRYnDrbAGw1FugCirfufK6R01OscghUskrmtyyYbAW/ks1A2G6rMD+
csevqLZ1y0k0WxC2e7TfrbtKJhZ8CBajyNtKvdNrQstZpJNLcEjR1GQTwpj2VAxo
4Vz61ZQhgkrgu63HZRQZ+/Vciy2TJuQyF7vpnfUwJ/J6kmJqbz0ICJD7JlHh+BoY
E00HpPN5puxc1Dm/EzVgvwXW/xruMic8t90vs/ORxhSOrB4XnUqHtp99dzI9KzL6
1DWmgspk+FPW1xVeKXCCnBtPLjGbqpymyPNuUdhZAVnHGhQWWBZXRq4YB1zydroH
ovMMmpcXO6NlZX23UVlV4m2723EMEVKnhXo+HOJy1rGyBvZsPr1WEA4C9ZXpXENc
UfV5aZGLaTbujqmU22AYGOz7QHYsFTbOOfDvmtnu/HbWuUQ1aDar32Xn5B9Clk7B
0GMn0SBo640O6aBbKnersdvuOSrxS0lgSgJb0Ht30c0Ts4EJZvZhkh63TB0i7ykP
oi5+lh0H1TcsAhA0YSxEsJjpUYxd+f4qPH8QJXKJPNIiJIBLXVVdhnNt4JobqJ/1
xpRuSsPfNBGfo33L0GVxyPOoUSAKF+i2xOpxdbrtSAzA1BTouWEqfwFqL8Jke6zp
ccB8A4Y0CwDNdpiGl4vrqyI4Kc3sR/dMI4+y8BbSQCGQzuUkmIfrW8yDD2MwrT+/
7MudbnKIb5Re5BlPTM857pSViSgseQzWWLLcjDO/yLMIeI/Um2HtsVuhNu4HMYyS
C/4bLw0SuGZ9VjujAJauGdMAUHoSj2XjRzAZ/WVPy7UcSox9zhfFOJp0BARbDeNe
uQU/Xi0Pdcr2oViFQ3UnFf1viovZ8YjA4GSNT1XDVZjUEkDQnyguNdeRIu5I6IlA
2MbiiPsU+jttLrkIWuF1hkeWVajCYAAEVNYd2NzxgbL0+hmoDu8I+bEadnxvoH6L
+xr5jXDu/SGOy0X1e927KAfLwFAjs86O1AKlIpLth2vXre/NoQVstdtQLemmtFa2
c+yBYOOeLdT5mDE/qz3TRQCW+n5x6ouXL2MFtrREwqnKfwnBoJ3Dr4G6wLMpBBvP
ILPUEE3npCUHZKUU0XrGv0z4Um8KAIKTvJIjL9Ab3/7YB+b1dALflYpItBQqXofq
pYdweTHmOvE60c3hR77b4X4S7B62AjYBmSXj6VoTSsBurCFMyF6KGcUfMnUj4dKa
EvuNyrdzmenSwgVsmh7ldblkhtELs7LbtEjPK+lKOLLka+3z5NWgNd7ORQfGEqpq
K+Xc+t/wqBznBgJo+U+xnQQV/2irHvRoUIWzRNiIEnvBJozz5KOHjEi+QAEuuhDy
bL3U+5aAzzqYTky4zLvQa6T5JzxmyTCj/Cw079DGAYPyT7SYvbi5mR+k/Hh+Jq+D
FiPxjfH8ZIdLQyY435jZeof+XdjE22aYegCfX6bJVaXrLm5N5OUpFGP6AhduOBrC
qNMOgXRJarDbMrQwz0GRSjmURH3ciuI2Czxb3NQ4MKGeGIgxu8uxPmk5sIIejAS5
IhwVUjyoz1eU82WmYiupvvCXvhkJAnM9d+hMDhPh0yrjrUFZNvntY7IoiyhEU0N5
MfOSRkU0xxYwezIP2yNJ3EU3zJGvbVu7UGvEbDtcz3IT3fOa3ax8MluJeyMsd0e5
hNV1QWYPKK67Gw30i8LrPjCt1rtVIKNbFU9hUR3ixtYP2uUXqy3Q/4m4H637HKyc
4vW6s3k8J9V5t8k+tRYmSokhc8bgUbSAxj7YQ48OfQf69Gm5el9Yh+u4GxZbeN9u
3+ToAE4+yWAIDf+pHRYgtoDFgkn9+XAneKxQ/6aONRZqDnTUsRYJipy2rfMMD9hK
N5cw5+9kgdrL/IJJ/LDltA+yXQWreCwUhW5nfh5HmXs/hiRXdvpBYwS74bKHL4ko
6X5rp8uNixRwFgN/bNJGAXK/X/kGiDep+eDA1+tGLB7SCX+v6tAvpwy/5qssLNOU
zr4OW2XMlww1C1Np5l1yc+gJ0QoqaFxWm5rUZbS4XstueP9qyu5kVXG90rDpG3gt
5JzZF4Cz5d32QaL3nAkrQv8OBqPv8bb0sRRVu1FMa/DRDY0wFwFT553hR7SV+zLX
AIQAtJpBzuzAmznVDEKg4q3o/Ru7wC/NbpQ+O1v+7qS3cl5RL5+uFLanJvxZeSPE
RWkqxRIX51Ri78TkvTWX3JY2FwmQEMaYRwGduQkglY5jd5T6x6SIrj+0IMlMHAd7
ysZ4TeWgKiUzyM01dtRaR25RRJIe3BbvCp98XxzJSuxCYBhrsu/xV3ts63xxjeB/
pnakb6F+IiZVIWFQPOT292P6CXHLUtQGmdATp8eM5ly/xrDLi+l5Rpjobrn1KzOF
YtPsCvURt2oJPdR4IajefRxQNbv7wJg5pq3bdcTUHAnmLS61bRjqYb173UdlycEF
GkQy+BCcsjerWINDzDk6lhtLZZXpGZ/nDy/EpemQiL2CgNmVwQ0xmABH8FgWjjh4
Y6QqpSxBjtUmrUSoEj4VS+DWB0AcPfPHSJWmw5e546aL1Rvt8pWWX8b89QNI2mh+
xZ7zCHn/rYAgBsx0pGw/i7GgLiO/d3IENmmKRmDBYCCN70bjAjhvw7laUCeJf/SF
amvKQC+KCZzsVA0eNU7PRjOZSIapyeolbbDZAjoAkMlC+kExUSh7huA9ZZqYi75p
fbhoSC9X4hTEOMZ0+taHzKAr+o5OzdGisHt+HVqGaL/Y193WFZTmDEdPa+GUJGcF
VBKxlfss85YP/e2vsg+nYnn8CCZOfe4K4hm78KUHDbdI7td/RM3GOYEZ3A72lY2g
/XyLHwjEmvb74JjtGr5GWFa9qexJITUPcd3ihyWR12lIKZWncsu5Rbt+wTOB7fwu
qQDyWxbRLA2QyLsqnzgd2OZ+M6OPoCoMyxq6ouW4MNCOZ46v0xGw+IrQ9Rzndgw4
bqoRIVMgvWv7aZwzFnmD2bQUGKi41CkU4vkmuOuz5+3BMG8Asr414wVJ7lH0kXhi
NSA1DSym4Ci/WSXY02SlRBZoKQCJ1JPiNYg+YXKP6ylDwX+K/XPyqmrZAhisAuWE
GO82L3PR1qzYyfiueyAxGqfaUpFLNduDjAFs8CgySYtFeQZjCz/PUEbQ9essiEzt
q3Thk32V+d/kgPoqVBFBXVU6fqCekTKkrDwLgblkPOm6SFqO7HRUKPzPYSSM0uqo
pRmK/1OEMwMNLAdscijruxcLOJ3lVtXRpqW3GnJQnR3bqPxuB1ImvdaouOAy6Hti
PFocdi2wiHplRVo67nD0wpOTXNfVst2ut3vBaJPa+Z7tG5vKNFOTdfb5zly8lDgb
KNB2IccFvUyaLl0sUWsuIA+pY6eE3HG+YA+GEzwf8FqOY4tNmp41qZFDsxZ9Esl6
kqvPXEaWiaAb4FugYoyQ8btHjHwPd42nw7EVHGviohd/0jDPJuEeFdR6RbGdBc12
pfNxyC3UFEIUPVbEibPAdHtdIo2NpPO/Sl/ZekYOiP0EvsueLKXJ8kF33Ocfzkvx
gArkBLO+qTSTN1rs06iZMJPnVPR4KPf3BHAftD2HzXKATK2iBuUwqjyu9Bj7aeNE
Z3h+qPV0pmG9sFsnn2CGnNhVnn5qFfs/+gntdUo48zfPLR9sSa5JQH0hzjL09tU8
aKWEzeu0yKJftFtgezF46+1xRKet7PutXpaGyQ7eOvT6lE324VTUYZQHuKgXDx5g
4voorbbKXXOrzDW+y/7HM3d978ZKUhlHVYA3rsHHoPK/7GEcMJMNjd05TXfMjaog
fUaUmnC3e1AufEt7MdBEcl/XSQwutc9lMBTpNzuwFLPObXy9C+yvvxbyKgXNGD0y
862R3xzpsmiZPTIpd9XlGr79xAhId0PwmQxqjrXX+8aDDU54TYnbzVHRwAhHcLE9
eXbZRvtAf18NDUO0zahkb2MyCX7Aa4cP4rBtMidqriU6eOPHKwDfvVGEj+C+PfN5
PEyr2tLG7aSBezShmh9kIDZXyF/qpGLs/svDfQ9vc1M7LODQ/z+pMnBdyPO49EH3
rbrEbJEy4WxAKWGrS0PLxlLaJsxomcSMKyzH0UGjCQjwiXwvvYgPZjyqBx6DdH0e
b38N8/4xrBciLF3pwG52BzjvEHaRlFdKx9tV6S6iDsI7trjWsvCiibRXlXb2t0zt
Xq9QxqXcrTzFWMnYOvQx+d2F5ESSOJnAZrUDwNpgtmvA5wVW7AsmegcY0epC4sMG
ClJcow1Y7mv8UP5Egfc0o0JjdZKYsyjXDWLy2M7n04tKaYI7whvSk5erXdLK/e5E
M2knVLdqJ61A5Qg20EuMYHPXYkCRw9y2pWQBpFa87nurbCZtTlSTRwDFP9EdqGD5
xk37dMP1G3reQh/139tyqLYQbJOBmQdm/qvh88oo5cmXrsaWsLz3OaJCjpVIAw44
NHmZdYwRTI2qUvfpLsPbZAjwGd/RXxfj5PBDRLk82VXCtpuAWu+gaFxsJ5nPZW8G
2VksJysN6pXK2/GwwkARuvAyFkRF86m/PzY5BnqjmBUR0Od6JN08Pjzf2ZQx5ec4
+KvUiisPrzVnV3VJXswYSoBh4uLJ3v+l0xNMXZhW+kYhpgpZtUFh91+DepW5PQPt
vMcpNJGsWTKMvO8ZE4u7+WS+LVegnr7vT4Rgm8Fxmg1dCm0psYgvn/4Tfo7nh5W4
IjTGc+so2eXs9XVoJpIcjyZD71YtRCJ5ISjpV7zDMRPHuRN2EBj+Y5bXMK8v3PW1
jjSrggVURROzJ+mz2NOpbr4mN+nGNZwWJQSXz6D1YVVTlcxjZoTEYk+vnepuYaAC
l9+llm5keY1wBqperZ4zZ9AMabXXQwJtQh9EJIH6lv5ol0jYubloJb+sU/AmyKV2
sUYAn1eDu9IcsW9Xuc8sLiYX+1VFlMkHZa9/jTkboqP5i1J0HBLmbZ2tEPtGOvzF
ZxuvbW697+01JnxNi22TgtwhwnerubR8TnmFjGWqDuJFhP/ao4bZZoKHMbsuRPgt
8o5bbHCRA1o1GKFUmEGIiTruMQ/9altyZUdfOfwX3pWfdQmAP5HFo4batl/JeCpx
TtlZjrSYwr7OxAnRRpyOntlYoKTA/dHluNIYgZ8qCmVLHesl6WnhUnUKwpNWY5Ig
Q/YdvhVQI+/E0uZMHo43vAn7J9mDOq7arZY/tXb3yaJKDpHGbdclKP7xxwfremFj
VvyRIPhMxz2YXOzgUCBRp9jrZ0uIc2Qm4npza39KxO10dvlICdRBQtH8sNcpAtZs
BjLdnlefgEnZcj079T/6Buf1aZQG9ba+6ILxOfR84z3X+YLHet5LYQDd9FsOerlD
qscxQtJGSPJE5DVW+58gLOK4nrCGoTjLZIa9qlS/vb7i431Vq1mfPUURBQ7OaaNY
Gi/GEWZr3qBZE+ob79TQxc91yS6leqhYxoPAbDeLAUAmsKOfRYPqvV+Q+juykdXZ
g81pzYyfwzl2bxhnL1X751f2MirKlHseLM+UzUQ5cRYZq95hRl2zUAd3c+/+IooN
/wnTWAq6L73Wf+5TNNK+aLzaRdR9WgOz8aCdI7+I1M5UvBgWmuuNgxNN2m6CzM2O
w6qbgJ7XJP1Wduq2VL6dAZ0sec060sYYTw6aZPuXupimHXDX2dGlKUVKfLjOhuMA
T/t6zu+zMuFoARP/Xn7inViWSkTi9njTLZ5bcLKLgSw2JMyAoFejKcCeoH0tyh3T
jW99PkqSZQCs3EKwHmg90FYDlCOh8ut158AuzRbIAZh2ph6SNEs5hSRzGyr2F9Pp
EMvTRUwLnOxW2gpW6cvDX6symmGTIwvyDwMNBbA/kJ7rkOp0OzK14sJ6ocNUU5p8
FiwTR+qHApHZ8wsISkJfSP9ZlSoBz3BGeFT5gnOAbtLFiUD2EPFMUyhqMZ3umqZ1
qVOTV9QUbB6LImWaPnBzBBv7zm+S2oB16l07c07XdzSMW9dPdhW2Hccj9ecWwBOp
Bm8rt6ZmdK+sYiQNUCEWm6jbYvu9stte/lVP8b5zAQubqfmbe14uYcr4rLn7H04D
3WiHXS+z8/ae6tb1mez/42+5alnc4pCLQfI6RC16KPKW4P6VEtC+JzvWhNCUSfJc
/ZUZrzop1X6mOIPFYh1S8EFNtGlypV27OsbUffO53HRS6EDHh/G45xKrEqN+KpXG
v8oxoZpirZKnmp8HpjyfMmJ+/buso3f56Rq90JXpT5vETmYNc26dSpVECfBSqxPh
wOrQOsDHT1d548keBJ1zgAKOc4zS+3D+xch2eX+mP29ep2O/bqPUNbulteFdvgMn
Kx7cSDHBdK4shSbge675QTv3bb3Z8f7c7N6QDtTcCRpIj3gy2OloAN5uWA2RO91/
DrXulngPhMguOZZ7DQyWyedVE3aaRgcZfXPa31bLIi1lHke7bzPskTje5c8QTkYC
wgIvRDfCDnIV09flrL/Est7XnGEW4I5i0JlkGwuFY2jJruAvANgJgfUPuPvFeB3c
rPXs9GL2S30YcFIOiomKI5pDi0qZw/h+o9kBzzjJwUPCeN9Z2arIVcjxctXJbwaF
NhljDxyMAw0Pkro0jMWpM5ZunA5BL+uXoMcWBNzLHzKghL6DrShAau3h4S34xKLQ
xKIT2E3mlM7vBTOOn8fkWcFYU95ZYBbdnx21+yTiUg8yXgnpErUtpbK1cPcyGZc4
5+68MSKa1tEACL7Hma/B4dnPCwrq6YoeM+YfspbIYJRkRAx3VVaNeABPs3zKQS3g
gbdiX4OXzLSeZzO+UQIMMTtmCC4IQsOLisK5v0Y/3zSG2A4HJlSUZtG4gjueKxz5
xZ/Gr3VOt0zlCCHs+2D2azSELmH5RVb+EIx4FqHVDYefJoGzyp9VlPXs6dGijwH5
pBcNz84wjZeHW2Y/rsFvL8F7Y4Ty6GBJmzlKYv0+ANUOPE+yUT27ypD+XzoPO7EC
1t3pQPACIQe9dywCMDZGJUHk4mrbKgYwonL3iSem54rReOYkwjuMPmzxcf39m3m9
j2THmGG53G+GHB8R/7zFz0XQRCqJJhJTJR3DM51/OlR6l9RQeNN73PbTiVuGzyIK
OV9DZ+FT/VJhcGRBSvZZvqpGUnPlc2DDysdP9RbCY2bLypWYmD3QGNsIG4P7rIE8
9B6zUyAuierQvPlg6bPGZfltjddtVDc7GSnEc0WQrzQHrCaRZPcoKgkgeL7kRAs1
j5S3GhJPRod0H3cAAiMdjddD66Z0UyCr7Xe99zs9m7i5ZQtiow3M7hgKH8MHny2c
kj3xHWYPc2P3O0a52Joe0sywjkFunIjA2yv7S9SvJUk9Xaaoq+U58ZS1AFtD+6xl
/KvwRbrKqmWLcSBCHY77VwxJvR3MekoIIjnPdYeYjGgoZIWoGxMOR6RTkV5dhIGT
Yam7/F4xdhKBL6at7E8atf+gHrB0HJD50jXdmGUp+buzsVLSwOAgBvAc+UsXyaaP
r8IIUeh0+lKDzSZh+G8tKKjIOASbquIEnzrpBh5LPFuAkGuOlRiJ7p4Gl6hoi2Ud
rqo1IaAr2Xh1my4tNKZzqQ2qNGUbwG/7quEzXaQy/f0XBk915/ADkF5iMLTWOas2
tqvf5Nc9gia9y91M7AazDwwc5sZVWP7yjcFnkjY8Y7SuQjaDSuZl87KmteaVTcNa
EKJ/WoLldI7L37HcWJhLKdNlSWKk02KTwlXySl6W0PPjS7gRFQZPQ8UrxCY5YwoR
HUhOgKrr2CXXWUE01gwq/5js3tzzwmcZO2IY7sdi9rnWIR1Igb2U0QZEoHYejv41
A6jxPafkvx4JVC4+icl3uxSwuopMnL8NGVHv6pEnQ93fVopi8Cf6G1WefFOBPgRf
e+FPFGLA386Oou0NOuTFsF1XBSjwymgBWCVrdawJqUxAvYh1IgcEMGD/M+55aA3C
YnxXRcEy5K0mfnc8JKz1gJ/Gt+8uS8az1ul/F25GcNeAT5Y6E00gFCucybAqCUVB
/O2Wnd6XtI2IzRE1KE6FiscQqODoEsyUsjp/QruQPyJ75m9JlpFkMG/RIWhuQ/1B
zdk9YM8bDk5pxmq9vorxO9FhPW9hSf90i4dszAApXAbiCb1qA1ywbKgCx5l8tMZy
ofQlndh7RQLEXiQUuEYs/7lvqq7yLPKyUgaQekuRAsK+lgdDjtSIfA70UGtg0pse
eE8NHNrtxnTqbgPp6A1y8ZkMDdW+Fvyi8AaE+wc6JxQaoa+X9N1TAB0dbpH4kpTh
qyEPacawJ7+slPgUMphrnCPyXY/LKgF8cM26FCfbxL/mjT1HmIqAvCWnkR7/Z8qf
XXZiZoSm+CbaZ6Sfhk0hx+CLBUmqY7/WN/5EGPDLPcdQSueePE2MXv750xBpE37v
roLpoZBpm4f7CvHNq4jV46tIebKcdl9kRSECRsEvkpFQM/bKjWpidNIIZbyUk7le
u6KtCcIX1im14aaglgc7zfNIfuG2iymcxjTLliTvo6nyHQ6JeBqCzoEdOjKK/yjG
Nk47LMKIRaBNYp0z+QF7Nm7AaWnfI4o8YIFT5KYNiE5dQHhAu5CmwXKw5H0GfyDj
7FEdfwaUQNiqNXqfJ2GhxdYTL4AK9xHIWFlJRwEngUxIJrpdZjbXRUsH8XDWbd4r
p/ZB87l6A4d5mT0kGPXeGozt6efs3GRz19GN+L8Eyx0K7+ROZ+tgO/4PQRhWNm4z
xAwjJQbjOqVq7zI90L3ZVpNeoDExD4aglnTpvvF58APrPGI5uAxrqii0e8ghLZDt
L4ydRaPe9N7IF43uqCWl2vtE87DLmgMBp7u5oDmek8Fmw/C3HRkfDnLsa42e56Bg
Camb03Q2znf81pXDTZVMz42o6BLyZ9U7lx/lmcEMTd1Bm/YEINv/7RYQhTCb/R9R
wwsyaINdYCIJjuk7LuUabqoJcmUF4w1ms0X1jTV5+5ffHXKScJQ4xitm5QLQGQ7W
bY80FeZxlJ6zy+PCLEAVefCZRX/YYjalb/OSAGp4Wzy/In43CDNlpiimxgPJxTYn
/zmhpetlfLJqAaaYDPHZHwG1yh2mnJrcPdFYJV9FxgDLaevp727OtdnHULrjV7FB
pLHODv42rAktgIZjeSuapyTsk1msU/Qs7szovc4bKEs5ct/ppV0TT49zrm/QXMtw
jOShFeBFpYMPYDb+Z5twNXcZtw5dQi5T6T2++NqWi2VYxrP+by87cXBHwZBVKHE9
km9gFO1IKxuNnlAG9BgOZU8eSWZWk6ehdSnVYLHjz3S8VfGHIuj+4as0kS35L99t
KW5dGRUau8aN76UrYFuJpZO8M/ng2PjiGTqZ6WvaSLHNcwyBoF1lO5jhOES2GYIW
3Uxo5u1E6w9LNyLP9SMWWJJOWK4DI/kRbZnwRJ553OSD/25nOX3dtvnFJ6hELLpU
r5ly25FAkjLZhhNM94k3Kngfp+7vYaH/74zKFU++LecvClbSZlYq/DaLqJHslbot
YDaW8EcXRyqAHxS8Ip4hxALpywLRkAuzM/65apRXtlkEqR9Ry6ARjQFOqaxoFeU5
v4vbIalbj9T0Oe++dNoC2k5wm4NC3AfWki/WP2R5Ck+K5GPoMU9MZh/C37ufums+
1qNBkXQFcY9/CNoISPAaiu5zwfJUAXF1MAmWBWrcn1QbvotgxuaNRRr84vXpyR6m
XOfFvm7YWD9q7to0uptX0X7YBgkGw9NDtF/RHigsLqFWkdYI/CwGgJbjsivU120h
d+hThjWCd0AgdoZe6FqQgPpi/jZ+/iU/tEx+GtY1pi3F2TqX3y8q7dfpQEIEPIue
6TCNs70D5lUQuc4VdJ3tZ4xe+/ep2ylR360SzV1ztG4pt9gw0i0jou62Z+QhzVZn
jiVOwIj6u1fBUnBwfHe1xEhFOIbCk61Xvsr4UDPLF/ihurI/MFnVBo97mQa9RDeR
fVfJJJ4ArEQhxZGG4MUKPFqrJ+vZk+d5+FYGh00gJAA6jqRkMPMF3lxAjXX7wKCs
5ua+f7d8xEUQfcWfFusgIdVsakwkS/HmMzg7eTXvdx0Dvr3YiOAKS9GfvqOMcGB0
JXAaiYdVBrPGWEKdnr4Gm0wnz+6Z/NEw9RMYJ/OBcIoPpeJMqrtv51gVjqCO9uax
Bz29VOTL8beD4/iFI+7dzK0aDSVm594alGiopQDWQiI87TRN4XW5Z3xLLgvA8jgL
w59VpbpRDXv52ugVi4ZNadDQvOYdma8gNXY1RBV7V2IdBUXrDZrFEkaykyzTgr93
vc18gl1A246gh4jsDWatUpIvP02b7dWMrI0neasrr/wfAstKd9F+J0QK371o13R6
tw0w0+1W08YKnTv/5ThP/tVFi4AEYbj2kXD5djBdFOKOIhA9drIfA6DfsnVcQAgB
k6Bh8NvlOs/K97Mx630wh/NIXtgXVNhM9QmXN6KmHJgbyPtj+vdmZWAnK3bUWEA4
3uI0JDWJH2oalGJgWC16OnxImls/3xla3oRMAwyFTIoQFnG3gohl1s1Ryi2sbDkr
MoLAXONgBiHE+9t9/qsuXN8ymWZec35fSeKMTZ5oCOesSH2T/YlV5m0o8HaFQVFu
+/q79rHGJBqFj330kzcTjyKOrXofoCiQMOY+rlcEMGJpPobBUvATeQznSLgIZJeP
83/e2Kr7Ex+wUQtnieCnHi5NP7h9MyvOm/vIBTt+8RzaOpSnCNzM54/QlrhW91Qn
Uwx+OnBbH9YDRvulDannhwSfpBlOc4WX7qze02uHtjCTh3Vm9aPxTnrZLGdwtC8f
I3e5UCSMxJgI7MqtjlxDa2RWigTmM7YviPEulxaIv2STXNaGsJHQkDvHpQIgep6m
JzhGfCHc7Prn8xStSa/6cr0+F0il4UvZor1pKnzT2WfvSyZ/Bc/xqM8CiepQGIsW
2nJ3APtaYMwiFFW7oZZRqNUE4izXPkOb0IytYPbp019hFfCcY2ghZX8S4dPWSwoe
sWRtEhAuEuFwtFbsJlZsp+RsDunboDcTQQVN8G0O5YTjrSE6ATUGivc9YI8YFK4j
ifJZ+7fm3yN5ptPRRSPe1kYrinrAIzFtTJaClgWND/IemlJuUCg0NHRg9KlnKnQx
uPfCMkf8QjLPMwXuVVUmk1ewYTc5Fxp9DJF6X0aWM4KgfAsmDeSW5nvM4tzHKYKW
joEwQC6VpGcolDnWq+B8KakG3OSRQvfidfrLB5cAPmcojtKT4/EKoWoG0RYhP9ok
wau0/bhQ06BEy54/dba0oteaMcI87N/1whiM5bzabbtqwM6kHpmZf+DAZs/tlyBN
GbyGrxopwVLaLYjwHcAjZU2gcfiUi1dBh3qrw4VLkF+b8bmxsPEPhcCtnq2rvzzS
Zcar+IGv1ia14QCqQVKgRk43fd9Fb9A5yUntzDMskfjIjSJA/6dlGB320Gx0qtcB
lmiHjttSL0gr9MrMFAsANGs0iDtkTRX/B40KLvIebdmpIAatcl+0L9lJ98aCIZsT
FsfRg4J+41DeCy8PlbizW3jCtMkZJHlzV0CTBALsrYbhMeDYE5UM8V1sFRe5xPyi
9PpJnH1JRCXc3IScugDcLm2XAim0t9yPFTvx1FSiiwXovBCAeRDPCBoDTZog2Ce8
FpPJ12t/uCL8CHZ6GMHW8A0QiD1GSY9+QP0BtIOBv2MOBVUM5cdIQYdgYsc5wfZk
qLLT5GZHsh6Kew7FDFqSxTtKglyDYRhJXqNsFAqTBO9p4X63yx9on1hIcSxV4SN+
I6kA/AaXZ0zMaRen8Utnbjw5QwkzowQxa5WB7o9bM9KnLbVzkoDb9qNBouvwux4w
4fYUakKHzr62YPcrAdp86znMC50Xm/rUmGwa6wWHuqmiBfP5r0ZnddMUSZms1Hjv
c0AvrnmVo1ywYP8q/FckKZfD4NWnm/TjsjOu9B5nwVO02Ztsxy2Ec83CbXmiRTwL
YOnFD6kgFhQEM6QtXEZ3U1r9vp9zH/+WiiWEzHLSgxOS8EUVMi1LMW9M4jK1/5Eb
3Sg8MLjVxDKTEQJmmhdYaA2EWgvpzy+xUcKS9MGX7hCdeYGJtMZ3di0WRs5LQ+En
UebDdaea2506jy8ViZEgjQ7v9u9EoWxbDHRdBrb5P/ZfvJWWdaiI0TPffu+PacU+
U/EsxpaJpG2bkcPMTTS3ok24P8lA61R3cFak5+iCkP7cMyBlkx2iPQYRXLMkbqGD
7eMEMZbVHKFZw066CdUDVr1eHUQl4gqrqE//nx9X9S5bIR9xccWMMroATioAPSyZ
FGJQDSy/+0PS+ko5sEEqr+KOUkqARRoplGHqere3d5Z+AslzAP/ZczT3cm4XcsA7
87S54RoJObVlZ8HjSrmCEKmIEN1Kudk0O8PGTJTZnX8=
`protect end_protected
