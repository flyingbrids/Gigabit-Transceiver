`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
cgvRlGVRFxoVWwL854gmrXtbehCaBjpt3vx08S0/+5+xaNT5rNws/C6ss2aU5EXn
Cq83IC64LmHm8v2AmfqepQC5HF9WiaylE1+Q5mpTmZxXbc2n1Aw5s1cQGq0deLqn
64/gQgfvMbQd3KuCyeJCwGjmzFzpMQGZGbbIOLJCBU0o4dgnhpZcxG4qSVp74zPv
9b26h2hPfxnk7kugfn23DTG/SlVK/qOwgC5t9JeIs3xPQBa9qJCmRyRdoWvXxyLV
hbHq9ZgcF9F8cgXqo2vQqGrK86Kkc4ldKJ43hu9Qmx2czhxFihhcHFFj7xqGj7qi
rS/6Ekpocd3bN3I7L52biA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
l/E0Oco0Pk07ze05xIrGuG5ivdRAtWpjjoCCE0wg7AyOGn1EvdTs7wP1v0zKJe6Z
XWXyAsEuQRAnfPCpmWbBUOvWR5jbtLm0+8ddZBn5lERIJD/K2egAnnOseVw0g+eT
Q4DkWGZfeXcMDH7nOkzx1JWuYGMNt0zfzYKvAphfMlE=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`protect data_block
9H37UI4joJ2EPokOiUDSHy2V84ZLiwyUPZlDjc+ghbLKa1eKMQfAH8JoPKkMv2v2
PrY7kTf0+KAejGdaJIKb4iuqMxQeLWNMJ9+f/G96JMEAaZpoo+FZjyQTwh9D8H/X
iNGJbWjeQjugM6gQax8jCCMEXf6GyW8sBWk1AyAaG4uJvwaHypMMFEqfXiFuoCgw
gufhVUREkegfgdFXuQTYpfhwCCERMYZkJj2mO1J9e96V6xL4Hx6RRbIjmwAbBMiP
BwC5tbMdTxmaSP2VkXuHa+n//S+Ms4b2fFm6OH7CEmyvntf9n0MbTa00AUUaOqCC
sRlLAoB8AfQITavi4hZwI5U7eMmqLS+szDIyTjmTx5j1SwoT0go8yIobBl6BHdRq
A5Vpt2Hsvaba+fgkhtH9a+eRqqPPt5VlpySYSvm72ea2LNZN56GSaGNGaVC7Fz0w
SHZ5TwDI49xgCig9d3a80VleoxgVcOPZeb1KCWll3JFmIImP6z5k3QvWX0L8LmBP
Sv1c4hyI8taaEtoBma/FQL97NnBvaOt10DnY/0IXrWyEQJE5/NuwP8S7CFj13Pd/
emRdMBW1nrXsb/zV9V2XpYGe9peXadUm7y3ZWeN94rAtAnvdfcmzq4sYtcd8p5tj
N3UXxrF5RrrXnlEyTVa3wHBsmlNkVRs2j0s952aXu1l2I6GJaYsuVwDmRh2h1odg
Wq20abu0Ak1Xz+aHxVD62+bK7F42uM6v/4sgTf0PVzquNRe4dk6QQnKcmmKzdE/J
vIS699Puef7dvnxtnQqQewY0QldFY9Z80txf84eccmwbXJvMgw2XtDUM1T6d7o+k
dweJ9SooIIWb2XXdPfdEfmcdnnNED8TZUAOd0c8nWcQfa7yM3BuXTZzzwDDEVWxd
2mB08qFJ/MD3+49vfx981D1U3Py24+mbZ37HIIrDOq6l2iHjMsOFaEu6yySysmX5
rT1Qa+WInruKmurq7aDf+9V23lcVwX+xIbXcEqaWvAIuGYnVqzivlFPGlodU/3gP
qF76kp24bEbPG08XvMCk1u7vH8wQl+xbfI1eLk/OX5+hM8a11fl9VbittBL0VLkC
sYD/+RSjKqd4QmHlSG4nKzO1WbiU6aL4ECUQN6b5B/v4k6rV6lnvmwFVDbN2bd4a
Uq+NKjICPbLpi1In71gnHRmmeDZUPl03XAf+vCk8nW2hzbe56gAStipwDIf8tnCb
XtVAxc0gUIDR47OHC2w5w9v0LI4q6WOwmAHLKDAtc8yjKsVa/uw9HY362sXin55E
ooXpwh5eCBf2Ej7kggOgEFXjR7MVvo+CS2ZbTVh1O2KKwz1DVDTBL8VwCHjB6A7x
htt3hKri5W3bX3rZDNd6KvWeNHVnjUljtCbmA4xOhWU56yzUKJP9QzT/4kFv7aR7
YwNpXbJTQjhKByh1K3AtEhp6dpaQ6UET4IXb/gdIYwsbesE0jdotM+RL2ClBtfU+
EKXjZqmlKkHJ2uVAHGi1Qg7e52MdOyzta8Tb/jGrYJdDeroYKXDNpE9JFRu9ND+v
B7TJ5CHQxfP9rRNYzuSCTn4mvS4L/Etjy0/FFB4AIWaewG4IWLtojRcqoIL+Pv1H
xzOXJS2OM613KfrqrXsYLDqC96a1AAtllhdy9rsXozKHgoLaMcEpkYRiYySUo8fV
K36M4nOz5EYjPSfk+ROcyzr3qKmElsY4Cwtd0pGHzAkesG/6JmE1HQX04GIz5ZVW
l6wWgDthVItikU9pHkhll4+gIJSNhUz099L0YDVwPZF/8HWwAwa5yXE08q4UNDjr
umoNrqKAkdwO/DPlsiqnSwWUpi3pS5CwBMxr60nyH07ljwvZxqY3F0pQqZ0k7DPk
42eBlKkD/e5iCdOTWAlpe/+UtYAB1hXv8G+EpfNVAZ8NFagWJqolOtM6AIzVAiCj
KRdFIRm8sz2E1I8h/mUsSIYJvGSlXnC4o2D6JcjS6iu2v+gVyi47El1UkdQg0YgW
ZZ9DJVBBbT88/zGgOnDPUPWkmrVSnc4ey1qIyjzQkzHvWBo9jSMTD7roRfTWnopx
1A4mKYdg728Ur5q1xOJ14kQBgMT2XYwNZex+vkXP6wMALP2DoDRXb6TKyUvME9M6
3jd8Y0a80yA0mM0lbnVi5j3+csJ3FEqa8oqg3Jxvw9soooUzsqXv7gzWw83TGGAw
Gg6RiueCr+1+5qv6Lfar4Pwe5jtnEu6ydEMrlj80uDMMjvYAiGR3dPQFdUKRUAje
nCHRLPMYbkCY3tcQoS3u1QzMx9mhuyLbvI29eQGl6xaF3mXKTcqUBfI7JuE5HRGv
DdvYPmRHE/itiUcAENtV/7DIUWm65c6aIlx2IfKvZtxgSBh+IKkkaaV7/qycl6Oe
Boz4Wz7LGICE40rw7T6cH7XrnFnAYavZaCET+WT8piHQfNXn5nDkqbjck41zHBY/
Tp/+aJxfAoTp4tWQPQwWqhmS1YJ9B2KO80MKNmUhCRIUzfs2jBWrLOnubYmiK9pt
boB3VFh5WabMd0r0vSzjpgnuyX/V+wjomJ/4674fCcse3D0TCJ4CQ39tnU+sOIMg
/s3DEtDa89cSOYT9VPm+bm28bUvTY71BzfQi9lXi+cGEGSM4Z/+uBBSUytgi1zsx
tDVv+W+ziLchive6GdJbk62xk0ebm7nHa2odHi+Rv1bsF90lB4dJK4IjHINO0wGY
l0iROEsittq0cqloKKMG64ZpEcyWt392fn5atuG0nCeT0FDUtjvY5DcKyFeoTC9I
s64lQLvnFQZ8iBedEar556ZdccWZJ/3b/Qkrv5Z60BJGV9kauSPsMqFknCdjqQ48
KRQGFup3o/F/uymjE819i4KR2DtsdaM2ygCKWoIBj/LK7I8LrCa3PC+QPPMRmwlV
2UjesX0DZrgslYBCfAPBdUmUWHyIK/u8UX5VP1PiTAivR/f3weqiCoGJJ8x2zuRS
E9hqCW67wy2WHE/ym51KYVGwmd4rccm7taBPidYUlygzguA9l1bl93zuLj2zZuch
AX0WlTOUlrxeoQGM/tT5QVl7Hb8xv/JYQv6u70AExZhev3X7UjFX1Bvae9Cbg1R4
QZrMW2bbbNgIECk9UkeOlreHpvjANmEotNjMVSCGZYwEKx2IYilILi7St//josyv
XTESq0RTvEBzptZ6yl+Oghrt/Hp4axZT5sdp50EU/il2BRCtahQeD13eWgHvp10x
g53vzmKJQx/UG2ycK/2fuJ0HgzAFACRohVG98m2ks/vWfZGzznzpZzb5benmTDWX
8zkXVzZhsUr8nfHlYBZilayF1rhmvJ/8OuthyF9dUDLCzmIT3zoyFOMFCdPpWPte
reTEjPu2U+zvQlkYe1gJdetoGi85VNhHWSWhFmtdh8jnH7oRw9OfBkEOriVh5oz6
4EZnqnQQTuqKcD56A5QOZ81A292g8qgfIurnhzK1hP7z7EyIr8Kkr1lnWlmTqoXg
Yk9SUIdRyCj7+coheQ/Ae3SjuFKY0rGaunD8pF2uO39JsIeBJhJx5kVkbc2qojJP
MbJXRNJ81KpGZhxjsbfE4GOCGFhvn3khRkLWaszFX4AX653DruiFnN1kW2Wt5OTt
bXXReRFfVnHAY7Tkn84bTM9M03lHHcqHlq8ZydzDT0jSLWqxq/kbkYTZhyrosrUL
3FrZSfi1oG3ReWasVA2z1NdI/sTyOK9tZMfO94Ge3ayq6F7NCU+JDxICc0P5eJ1A
ob0gKmq+aS6RB/KCnznQE5gzCRvBdWxEYzGYy7jHlwJDNR4H0dACPGOL0X3OoxNr
dGYywvgpnE2eSn4+5r/DsHHguc06AzeB0oBpERUHwUhCjhMMq0Y2UzDuxLzVZuIO
UobtHdz7Ax4zzOsKQOkQQg+ef3EFbJJzxHun05YwXGIZk7+MapG8mqMoLLE1TOAE
q9NVLJJm9QLhFpwdmVYh2IcDog+VsB2nDTTIf8fD2ijB+1AaCEgQI0xMMiIgi9fe
FxW/mN7+fsC6Aqz421qADw/jHFeKsULpPwIyRgDAzwNahYjdDtH1Y6cZZWgv4ugp
lUGMiPh7Or1RnpuQPQHPidupUrP9wTRB/mnLK6Vh4asWdBLr1Q1hfkHzq5HoBY3L
hPXxuScEgOkYuv1OCEO8xihR4XoIkSlJttt28CDEE3f1TogtFh6a7eAApbTQ3Za7
lbaobXHyqIgHm932LdB5PT0qgg8c4l1o5eVsebHqxlZmo8k4np8bFi/sRGGu5vSe
WM3BbVxvoBZHxZtdd2O9QFb+KIRiOxewXfORIdPi1gYPC615xl6lVqIjmI43cPWY
mlnYMVlvmBCr+bLnHz4v7Ici4qZqyncVyQ86vsUSZ9fqCfedlmMNBn58/9UudlXy
CDrWwVf0rcRcHgbWxMveIXiUz74E51won15lUMJ4QDMEZvGbSS+veIPRVQbRrKk6
XENTDB1jvKURmNmZhaTPB4Ffw8BhCbUGBco5rFOTWcVALX5dkhql2wZeIkgOVlHM
YibQj7ILoMaafIK811Wv39zEA/VHPBhCdpsGLdZYdjleaEhNnFyW3y4IhnK2aPwe
ITka2zm4O+81WMz0Xf7AUIEchatPXoXWHELA+IYt5hGP8aN1dxCDJsVcns5ExvQg
z1lME/U6FNR8aFHKSOTMLWX6f5yxJSU9tNB5f+hZ+wgj0cqjqE44NcNQ9AVhSLyf
IqB08GTcVIyqIU6XygAeLbp/jNmiQ3hiQfIPc0inR6kS7bzbMzvCdALzQrp8FWi+
Rv4bkaVzF8wYMOyrRAkb/HVL2XrA3KG5uColzSPoYVOquomRuxmUFxSiu4DPztAa
2kSiimGNIiUGRrvmSuzlQpiQu2kw6CS2lqwhSM0yugTvnsbtoE5RQibfkafEKxCt
LQH877nfeUDsQL3V1+tdr4Sh+xiwI20Wt+hFJPwGNeJGBvyaPc6KaRQNF+OQ61e/
jmB38bwXt3zzgTt9QhnBB/ZQ3JsXdieLtuQy8i77f+Kfm78Vj/R03jSHugRCu9/W
1wcij2DFjHT6xNUxQq89nm99uKU3bYgUMj6Jkc7C97e836KjI+ioCZTb21GGumxF
oiegaxL/1+hhCxQqOv8uQ3+60TybFTt2BjpZsf2hNi50IwE5y9EbF7CNy47TLaLf
Bxuowdm7vxPpzQY5OUQV8sS4FUotgUN1FUi0Hdasc8dnEaFPnPUjWUrMuCBv5CKk
nSmXQyTEj/gg75qe52EJAdwzuf47gU55VaBaU5OSfTEdX2KzqFjUKmlezyf1adGI
AlI5Nc+VEXzf58OBBGXVJiL2nrutPziySimrGscK84CXPfcrMVgFuru4oYsXaWZ2
NWptLQbAEMWySpVn4UhNMqF+kJPLxFatvBXCSSYdIw3SSGEvkGCEMUPyeIS1AFcy
mrxvaZ286TgYKXQMcQ/ZizBffj1KAYz2TicnyJZXDzMoZSIw82mVpCG1Zi8h1GXG
O1uf2Vy/Kr8K9xiVOsFbhx/6XJksVJuyw+EZ2o96UFA75JtsC3lCl0RWxFYAuqUU
LSVKsfHW+VnB7Ujn5Xk6M/d5bnoCKWVEWToJlyxwHEvhxjgpm4WM8YiKBXP+oyEp
O5zBrBTBzOEO0bgUvVL7L9wXTY/dcPKwZcBm5xSHRA/G1Xth8t0yQrxCOwB1ZqmW
Z9/ndTnbzHSXrnoRyj5LLWT/ihcPcZEQCKkC67S3BF3pbTsQ0nbziM0AfFGeGqAe
6h71brRWntGZ7pGEeHdt4k94imrSEfsCvKuhronSAHoPbn+19XPd09v9V53sOi4G
8JfwhQ1fk8zN1pXaw2y0Tfxhx1AgFkhE8rvsuuBfAjokkcceBT9HThe/XvHTLfCK
IO4lz9Te7pbxJFMCNJUPFaXZwzeIytSigc1WqmRIqRLn7mPUNIVOlbG9h87rQ+IB
iQ2zrAeMdft7bxuLp+1c38oEJXdo0Ujn8sNwQvEKUycJUyhlLFjdNRzj/xnxNRAR
qGgsVk2BX1VF9qoHMDy4GuT1r5fn3zrdOB1aeMgFsnF/c79ju8nS28RhpKaa/Z7z
ezRi6Zvpc47tbYiiUVceCRbMgtvj1Mc3L9cawHdVHJu3ufsp2f0hcOv/5AyyDLhF
PGX0HHEbbM7mVPgIZnS8ztKkdO+Txvr49wxX/YdGuYxxRsrD6QeD9C+acWaIm/TL
QsOnnYZQbGT9q6ynqotvh5CKHU1i2+xijyOCVnb4KbWzyPOPCO1Uvdsm7Wf2ZqCt
KFZKj53WqJ7ywsBfLbRpXczH9t2zFmXlNFtTTu6HzrrCqhLRbIr+hDjTbZJf8lhF
Enp6TUe36S23DNibF0/qJlL7gfbbvbxHuD/akgp3rUO1FGv46DHUJrJFWPS+Spno
lgi3ux1CpbK8qwoQX6dC5/AY8Je/TR66WSevDLST76m2rONlZZHUsaGOcMLsVPwh
8qdjIy/nhNreVZw/eSPn6OOJwoaeaMwENxe59nftEzqHbTNiBTAymVGd04DID71w
NgAxbcu4R0fIDJXxpR10AQYMtUvHgdFmEs/8lXHSJAeg25d48EBlyOONm8omypPC
/x6W0QUlLu6dI1MiQ9iJdDtAAGUZh7Ui/owqCi+M7fCDD4Chf8jIvzUdAV+kPLWX
b56T1y0Zfw5SXzWVZxrEqRE4A50OTLnBwVl9i6rkpxxhzQB8VA3T3gFqigJg32Vb
884C8AZdVMrgBAGs4MM+9ReDjCksSaRECIZQIIVYoM/+NJAzoQYfujA/LyxHobQX
vvxVvYyjD21qSJ2z18q6rtfWa41Y4cqDtZDH1d1YfPaJYUF7yEYX3Nwk81OKpPx/
M8yteQlTjiILdiKYaWrCt1dZNTunX9+nd084lYZWbA/qwioi9i1FIC+1u2Vt+Mic
NdWzaewW9hvvcL8mDIcgsDl3YB5fXXwTEAg4X6GOOTVaVwwMjMxBOkON/0MXwpdF
jRrgH6oIndGVTC7dAEWCXWjLRd7fI3uAt0rT5ph4RgTqVWrZlmSmXC5WAu4Kfnbw
6UWq3RqHt6MI6eP/vSojb8ZkstF+2g+9OS9FOdwJCx9bEltSwv1HsUep1RdHq6ZG
0b1HxNHDGFBEwJs23ZDtfaOoc38A8sPrmIYkF0EyYdsEZNF1BBYrAuBt2Hxud26x
fguBIW1P4W+XRVLERZk93ORvf253FtEwPxY4HQ4BVrxl+OfmcGMzi3BFizKftKa0
cPJ2C9P+8FWdhkjWl/rc1B85Y6OXimM7WDJvv8GEgGlpfWFsLA3UBJHeatMvNMcS
D5bQJhTnap0RrvAjSlsftcM3a1ddSVVG5UWWCAg1NWzSDIYPNQY8fufO9pBwq/1h
8bRT7Vg6JmpalmB7R9L/HMDmRLaX6U+4vhkqm+5uaQecSISvc/LPnYJrgNLf5Ri6
86GufTXCsHjHiybji6WFIN8YImlQCWQopBS6eavWGxfzzq43Y+4WHaAbJ9ph3qam
2Sr8pPB6L6d2N+IvMhfqWsOuarbPoaVVMONbRHPeWiqRjFLHikweLZK362BY+v6d
zLWABfV2ohrtKT38iHX1MDEDqd0oUhjpC3+UAwL3qy5f0IRkygghYmzei5Lq1Km8
`protect end_protected
