`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
N7HktHTrwL6LzVjOcJRmLPIWuAqRSq91mQnw5yz8iOAWYp8/33adwJuVzd21SkfM
1cJKWnflHTlDIeZngbStzFm560vyj6uq1asxD1KrIZ+JYaiqdS6dNB3PDrLVsnHt
rJvyhQ5Lb/KrkM3yQ5MvMDZhgInpDWOZKM9fVjKAOz5Okzs17q60jBrp2fJxi5bN
RA6co1yu7smk9admUf6jWBWXo0o28eQ5DdFbr9qnK7Zebegc3HGf48BdjzE/JMD/
2zcsxlsfFiEAEZGSt+fpk24omUkZj53lpDnubyzvrHlbWdzRbESqSZ946TKyCXZ1
Q0EDf5w4j6ZjaplKR6Vo3A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
G1whrt6iEGpqIsFhzD7f1r29x9Ft6ZDu62y4+DiXqTEEGrMLhXoBPXFu5j9hrIcG
Kj0LjIcWEtGM4oSpbaa0c5LP8HDYs9KpCNgFk35XdhV3PyWYIxDS1smSGvx0nOHw
tR9TRu+x3f0qMB6pgbAe0Il/mDTldG69JH+vKgy0JcQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15504 )
`protect data_block
gfydnHTxNlCXNL4qot2IH8XpvwALPnBB1zrAdY1yj0dDtJ6nFTPal77KITmf1YEJ
/ROLZZC74IBP46XnfXFzAaXsIXOsPdaEqkuUSgDrVc9z89aqndR4KVHTtkt91NXG
oK44xmCQmG8ak1awbCAyX+yk4Ni6KByfutCHD7YKb28OoL0SaL8YkqDTqLDKldk5
t7dN3S3WVcXtxucZcKkukQf3BIVdWv34gSOyPzK7sTBLMIA8Pqnaj3o/K4Irjsa6
JLRoqZO57r9YfN+vLBnzw2YxwoFKGN9kog9AUBRou1Ds8FDIIYDgScAYa6YDOqWU
Mm5DhS6XFSnnOIUjlsk0s4R6XwYlS79Iz0nNcPZp/xIzCS1bgnml6Qir63nJ91tj
IwCnP+ZAjy4X6VSGMq9IAv4mm1chZ3qQ/WPCq0as86plXEjSW2B96g9kfoDA9G7R
22SoxnhrxyqE8rSqR0XlGlf+GLAmCoh9d+w6MbW2u0pwW910jjFCS1VHZJMYz7PH
ABTm4QkHyF0pMSu2+n+L8G6oAjwPod0ITyEGDctyuhK3lRz32/ef16ZjsnO4oCkv
8xI+wO6u16h/14hJNOZeMbJnlzxow3/6E5hCIx1vtR7mUIWYC+TdPe4oiXPfzJqZ
5OGvsw47NjreyJ0tYjhKJaYEbO4X7sRPK4g9qrf28FUXMJs5Od8V0a1WlwYTwj/T
QQ1F1fYbHTDDt2LhxzNpJ5RXitgL/0uwsHDRJSLFcP4czCJnnXXGT2DkI9o3B8oy
WAHvLX1gDhzYYLPrP1UmeLuoNfDyO9E4fpJwrz9QkiUZFIqDT3MjxmwgJOpyHtrt
INjEB27OSmAqMF0p63Vzdntv/GULo8l6PrLpyhKzTlW45DVNDuTJMgrX9JAYkolt
4SS6HPXFbiZt7RcloZUV/ZUGth6ppDYjHnovNFGumXKbc7cej12GZXax9wyyFdUj
aK76w3I8GkYvFXptQ8gv9BHxCfcu4UX4Vgl8VWm6ZG7ZQZSkHA/BMiNP69yFB5Fr
9o0rqGXKoWvUrdBB4FA1TdAV52xWeQ5nnTetbu0+1PeZZbr5WnF5kddCgiF5YF5i
ptSAYff9PQmCz6WRngHTUpGunxSZa6NhCowa5MME3YPgS4R4eia11x6HnQcamDjp
2XHzgVoDhEjAGUC2Fyr4Xd4ctgJIBQ0AZkbE5O8Jfja56cGk8GBuWs6UfqjCKK2x
RPKPAtlKVi6n2Mr9TKhS/rvbH8py2URMOM6hWVlInG8VdTNJwrl3zwnI7evMjY0D
VfOOV0NGaJQsh5OulnrS/a6jIrhc9hIYSWFTIh/L/eLY4kYQaniRk65D+NK081iM
h+AYFAeZlWqKNqHUvCcxVEStguW33hWMc3zroIrb6X5Sq7/W1WKdbd7HfbJSX+Zb
68yLr2wCUeJXIZtY1IhtQV3gmakFMv2xUq0z0e0aki8Qpg/xRukikfSQRLcVtrGn
HCI+fj8zth1hYMz/59Eb9pCTqGICMGAy5PBqD+FaqwOw95M1rbqwUIu5uPH1vxf3
3FMYWtzdajlx9v1l0qYlqtzANX7z33IF5vrtSHs8xrJuie7Hds+crpxtFKt6nEIs
jW5n0zxdi1Almg/uTRijYYAQVk7j+g4QincmQy0xBFbk6Yb/rNw6lZvrc978WERN
JgvFrlLV5N5oWk11TzhNsEWMSNYIlE1Sv5dp2ES65J5jwzNhghr6bWMInSsEEnim
CcsE/sq2rAvcL5hj4QEbXn80NTaVFq1hB9UvGh59bdxSPijCQLL52GWqx4wBix8K
HktASFXDyC8s1IIr2UJKn8rfuXX0HJ7vlxKZjoLlrTQOFAVytjJdWDpOrkIcfphV
irDBhBMwrHiMk5h4wxb7C7mg5fDL1zx55JVfGxsjLee2xE8CwsozR7RMcDFkb/ks
cHIZVb3X7Q1+R7j2FEzX/3PrAo06TzeXYKoiDQn06QWJcV6dw4TeiRccivsYfcCO
t4uHjgDauQx1ou6fm9Bjb6rvjRhZVPnwwDLG4r9FPwuhgiVSpGKg5zFPwnL8oxSZ
AF7hluC0ajf0aDQ4NOJfd91llFwRgp/U0XIvBW6KjHiJsx4MWtSQrJ6rK2bFo04m
fDlskbX4CGw1F6eT0210w99zNLPOWQR+BS8TALCg/u3tr0BpXmAV4fagmtF8KO4R
BPK8M4UXlrIhPr33dM5IVi0L2W0uPJIkmFfHOkbrYYO2iUtW34dqEJx2bvNboVtk
7ax5MhxrsOfC2DltwkTTN1qevioMUv22LMc+Ne6/Ld+r07S0xkqwzQzaM8c8IKt3
qDAFvTaZNroJ4dOqglt0SL523rdYa6gHReDwihRNtrUephWFVlKceQsriPrpGH29
IPGkhIZfymLjQg5SkmPsfrFe6BVkzH0Q47jWVeZpve8KxHURCER4ZIA20sis38KE
yeL5JhQlOsOkJQRt0Hwj5UhG8/ihhscUwnHk+uh2/Wp8s1Tv0Yv7lZy72HuPkPB2
KwC1Yr12qPuCNNjqpd6DGFMeifIA6L4yS7mGxrqfoDMYLo0t9WW1jEvT6Yx6t66O
K7Gxyasph/twQ93MmMDXe1wge7k2lbeLW0i5WL4IW5xIx4LnSEMlsyb7Ja+VTgqu
3iHV7KWp6zDlV2n85k/wtGHYeo7DaFAJf7WiAmgvgwCvgcd4IulScfyyVObowiQ5
t7NaUVzNhkvklGw41PeGD4F8/9kWCMqX5b0JPFjw4//MCbFZKUO9aMXNdIJaawve
5R9e1dISknojWZjfYs3FTyCWXHqaqWXp4+6FzRQjsA8Z/Q8vMuiWcUIJPLw9rlRf
0WcVkNB23sMWMxgFasZCO3TE910YqNJs1T3PUlWrGH7J8TeJ+jzA0kOzZc91nVm4
wqGlhJVK5cBzN0jlBuRQKVtonkcXM2v02RUxIPy3YX7+bBzJBNnJdbmIXKrmBwII
KCPYWouoqH4Z9lmQUPBDYEB2ujBgO6SveXj2bqvCdMybCBEjs5UzqdTBMCOPLjlv
eCqHbuet0wwK7APnE/gRUccaoWH7j92Ii0k9OXj3R7sDExFLsHmcBimBhS8oqSUK
AZPyFklF8lYfS3k3NbkWQiq/lK8h/Ka9eaIIu/1C97ui8lQv8s//vVgOEvXE2lPD
eEMyoBcit8l7/TDsfqlPMMgTEZOCmSZjAHO0BHNcxNMiugfB1RNqRE2TxwU0YCWU
C2LlsyG5OlvFSmk+JtuSEqaSkJABXcq5Udj3Wj0QsWDDM8UT/5IT+DXZMKRCGEhG
XdHtKevoE2HJacacP0P4gH6k663pPnBnGULe8pQA5b4A+mU6hzB49YvW5K/h9NvH
VL31kfwWv7+HKBcx4E/SYkTrjIQamPrx8t9iXk2gvbS3mZy/VVsYG+WwFAto+11N
xcD3Q2dMrQTYhKrlXtaGGpwgyP55Gujgh43RxuBryfKnbCi+3SvMPO3iDeSQ4Wya
fGKEpKSa1z74132bFv+q6R4zd9VFn1Hq54Nl2KOoghEeojRQYXtWPZRljvkWCkWz
Oq2r1Sl4zhD+kLGILJTd7cfjwgUuhbeUQjSxWU3+2SQrGpqeKQaFxSAaddfVD8zq
NiqE1fqSjtQX0/F1eqj/cm/tOLVemQGWd+bZAOiKB0V+Jw4gAiu/UV5zqUPL0aJp
hQSvRluDFcidJf1x8XSCCuoS9bleIxITIoJ2hnQRrtVyjENOmu7gXcEkx4OtaP+z
8Dxrjf6jzZ4ZJcCoAWlUFLrwah8MnbsImcDkAX1iDIhOUalS6sUX3ntINIBPieTy
4J8N+lnyPj21ByQfhlHheeRXgmyEPspyqPmc2oMsQdp5sBj/Sc94aDD2zLiGrDXE
HHaucyTOBg9Tg+XbmbSQJJ4/5oQ+QT1piK2I3/RtFHGBncXIn+DMEPYF07fPrYAx
xepz/ogyul1r2Sb3JeI4vJv6JqkxB5Jvwz2F9DQkxYbTaULU/lwUZpZfDmWBMwn4
kh+YgAqtlsjb86iW+VLB2Ath5n9oDwvvaOdvZVJ64KaTOEoiy8Kbo7QNZTEW5V/u
qrdZUejsQAFZ+7Lq54puY1cGsUCc5ovOkhbA11NIt4qPSjovj1XOKxDMRTU6zm8G
VrcrtBWOjenD1YwSozF4/RT6EUi8Z4Lu1i6G61VknUSz7hU9GVVqzMz2jkp42Sg3
4cUegakkQmTwHafzNGFga41qeFuGek8yYekZ99s2rARntvzuikt80yWuNs+0mP46
m+se9XHn+RDbtrO92oDzfriN4+aSu9CZG+bRe1Er2ThvIBhT3Q7mO/1uveaXhoaQ
j5k58vQfLsTBvNzh37tMByxy9aHKtgXQNzEjsaGn45LJsnE8TPiXGhI3SP6hs5RB
lPM47GB/s/Zqgh39ZPrzLnA1LtqJxQn6va0ANyoqzXFVhBM+V7pj8+0c54IhpR4L
20rLoyt5xZtO0OUHoK0fTg1IC7JawZs9Xtid6TcODMLFpAv+bIx1XWT+Woy4+gFu
kJ1jnA3qZqb2drH0hHojznULOofhpwgrK1TCB0JV0BOOEk9dZVgodNGAgSp1oubV
XnP+7k5VpzYKFobd3JmzqEgmOMINNgo7pbcK44G1cFtdFLwA8wxH+8P7aOrjGBtz
uEpWYO2NTcqMsxBTfIZGpnsyOLhNDxj1d/neR3xjuzGH9zTF9E5Ixoz8PYEQZsyW
TU3tthh9iQNdixC6G3BlCwtVYhPIxR8FNcv+GmSSeloAuqHpvEBdbSphac95VAf8
I3hH4wklVR9aIXMBGYuOdCoIjzUauCbzVFhQRFknNmWBuLNasLWnM60o4/Ul/5pe
iYcB+De2sWELBVg/FUyfM3jnBdsB/5yzUtNjP3FTrOL1WSwZmKd6XnCT3yTHrAG7
NccNVIvUe31l+Gu/JkNNLuxoLdDlyCX+7TANK4N6lWod2A82zBIiAvQENZ83SADQ
Uux7snhOF1IIRNEIwCtDyf0YWvYFpVzAiQPO9mNZ7pcIl4FnOlHVjard2egkrF0I
TLKJkGs7gtDUFSAZ1pNloXWbqjIQIHwQoqMgkRdKk9QILpxNWjf+2UIlYEJWgn3I
td9vIvOJNwT/Fy4KfL8nZU2J2LH1BmBDR4bJpgUKIKMv/2G3AjHyLPzM14FUk9x4
/9ZjsJFH3L1/oo4AJQkowNYxCgIJ1JENuBFbPz+5cUlI7nBR5E+dKgg6vlldPJyh
H8PD9H/LqWb2BqQBrpQD1IbknRP/e/YqcpeYooaZEUVhxxRIa6zIuu66po+fCCA3
7hU6ufxiVncHw0OE5fi93+ZxKt+AbfyYwIHHa4sjbDzOv4dPWWMccEJWf/9MIobi
2aYmpcBWz+yGn0wnrXp0kS1A7YnYBxo0uda1ugcIpCL9eJmMPpOtwc/UWvzgGolz
Cd8g6sqee06H153B9y+2YDr8mkRa+FfQwXF1xnN75vBkOII5tSAufD4HBjVz+jf+
eqMinBATL53m5hkj6/Z3PW4y5xm5+NmTI04QmXSvVzratvUY0dB7wGWy9dyo1grF
tMP6DalFDXICTtgg2dQ+IZ9nDtASgeAwb73RDVbCx8WIX0FdOQmYL04PQ/KmF1LM
v49vpJ1mVzSlaxvhcRO8M7VbcYs0OlwjwvWYX0zzwZIyy6xKGDFaLtxfVmOploRd
az8BWsYLALu+xAQpy4uo76tF+rgnXKzQgNEReLOgxvRr0+fdTOhp/cK2ORpe9FYh
/KVNG+GzNlDTb/E9BdpMY7HU+XYjIYgb6YPNGbNxxjauZqoTtkqsgYmQ7U40jTCZ
wSbtlgQfA0j3hGQovTPKTD26+yMnYzumE3u9wDUY7ilgyHQ3KMweS7GntHvgTWoY
vACWMCI53oFTfqwEbqRaP0YHNA5GQj3uuR3a/kQZ9ezvlzFcXlmv6xeULttuahi4
xekUHRwyZEFQaw1+i9hpLTyo0XBaqWO6FRdwLfswmVD09L3yJC40sAqvpV67L/8O
d9k87jQCsO43Q8Trv2BPWn32walZ1X42f15ol0fsxg9KsmqfUPuK3UUlP1cyzkQt
Q5s3lP7t+3ylgXJTC1DULzmQRj7ASDWIaAn48y9rGi5TeCI/qVB8F79QBhRl5GAV
2+WJimq3T/xWsF0nRq1ZGBj9Tmguv7vJRRKSPTPBpfTKfT40p8j58NlZywWFy9+o
kmU6zL9JN2YOklYW8sELVNv3yuMykFqMAJ08ITzbRVLpmsWLUc5EXxhKwJi04DqL
1cdsEk1GLUpOE8f6WCSnm2yZVXc+StCZDY5L6q756BMu3gXTCX+nZM9CryNIPx+V
VPFgzJCHFSBJGGGC2QfmuuW6C4AgZgSspdxiRA7NxTTJU3wUDMEFRkYzh/kF4HQO
Huc6/r359ZReXTzMruMXN6fOPmw9c9t9KWrYdL+yL8cTAiUdP6pb+/D6zfOIzaxM
91r5kVW5QlQsX0D+232bDHaeMYVHyG+Ws/FrP4HOyTuvJwINIKG+RBI0X5KBzHpJ
TpzS554nvMa7nyuJXsCrnKtwuC1ce91vcD28Ego9K8OyJT0UhH2LWtEdUekzJySQ
ggAhDCNRPLVyWy4//B1sGU72qFvC3RUBNZ/UHTseFVqB1Zsg6B4MPPm9RPsDGTp2
5bWk5EQea5Z49znS+Vy12D7G6R7Ja81rQUcFYpFoOHVJykticP2xFtKpY1WSYqv8
dzxX+wsCT9MpMvOyGZY7dH526rZeMBxRg8MN7L48g7L+zq2OX1X3DNzeURvGEMdV
6WsNUxXrFPLjVmVXOUUdawDlLqW0z0jFfuC0N5N8W1KfnlYOLndbVaRJ0/JgSuDU
zNCvwLTNod+85v+gbIPGyMM93r6FXyVdJvbSUkmc8x6cpmRhFkQE3u90WdygpJrx
6hRTSfJofrn05k/8mhyu2PX7msoPocXUJUnsYGpqKGQTBa+YfRgsHnTlVMUoe+oA
lyzRqZPdFFZY73l4pPiV8E2/zyAHltYQxp5Bg3+vENrnQZY6g+nqhqMrXt8wG2pl
2KabAd33xtTHTmwPEp8kE0xeWXxEekTbWn724qeNmcqWW4T1SG7ZFOsnpz3IbVHA
ikfxnbGZRmGh43wrLhK0YRwxkb33rucxaFHdfhgaSI96EPH3V1Bpq/2kUC8oIGul
b6Lc/ZdV08FcAAib00iMUV+MxyaSKqrqIgzviPkbpVV59jr6GFC+bztZ65dPbrOa
6h2QPsurDF2miKW77eYdeTjMucYiwwCEM+qZgiUwwiCZZ7iu5lXsu6CY+M2+LPmn
hvpRu+L5EYVFNyuJmNEErjufOxxPAQrMkySdd11p+iEhPWQCqXUS+TFfsaPTo1iV
GZtRuL0IPj2yzVio2zlQmNACl3rla1huSjbvCtOJ4elKu19kLv00XbTYvKS8RZw6
ITos+DPmlNmOLduwxPzGm1iz1CF01372C4EleMLm5pdRlpTVcsDX6McGduJmqJBt
+7Covz757YgLYvb12sxvvrjOFME9P2wjDXKLVyEIy3fxBMKtL5EIbVvmjeVknnBa
+gSi+e4xzxudIAjOxcTOK/tfxBPzZRXk2wJZheG6smb5h4Rq26zoOl3HTQapErBq
n0tzmdWrk7AozomBP0JXOLIruQ2D5VXSb7OUOkzz49kqKPgkCojdEiFvIOKFddw+
xmDpxokwKEoMbQpFRSaTiuypE+rp1KRe+SF9aRP3+wQyKHeDWqq0ZVkDG3yps8m9
ZnUgamUuN18383j2kb9HeNVPnSQs4cBo/axbhsO3sirvkq2O5jqOF2MoXWeDmL9Y
GE8SRf1WvEO5JjSSM6Zigzl0Fkk0Ut3KZe4fU3ev8zLyih1PCxzXEpIvwvX+rDXc
QsDBBsiPy3s6zpYszlJ1H6+6nlKmnWkd4kCzg0dggbgvHXoNgFVq5gb93uzqY/jJ
gSj3eJchDB7J5JyIyT1bQLE9gdUnCwROOVwnH7o4VCqNmJwA17aElMwur2oFjNku
rLw/BH1807s0dpe89d7z3SACFnr5RaRTdU2ZJaX9FG6vf6uM6RDKCR4h/X3LJtAE
UkG/Aejr42pn5PmJqT7zV8m56ra+PAcV8TstzbGv9PoMgfG1VBEscmYdFngmiJ0S
q8io7ic4b1fF7cH/FDduwnUn5zqSgUVxtfDDmGP7Ju5VWKfvIfKxQcRm5vWRyJFz
o6QyVX919x6AHQ51P66G6uxNMS/4rT5AadU+10a8ViNs1LYMZYvZ6xYM5rtqEmYa
n41ogv9H+sYVBNaPhwtvgcIEgTgTIj06u6YNHAP3bXN8z2QGHb2xWHEys27aSuuB
3BSwR7ue463ALI8bKmiwvuRy437M5hp8M8t7Ayo3VrSGTsznXnvAQ6t9oXZY92ud
pI5ICjGLRPLKImxR00apBPBPwi3Q1QmAtiCj/HHNfcldecqZUTMfAyNyO6tL7X6C
heS7AiT8kddR5oCosulJho0Od3uQeaDlCHUNXcWGpCvJudOFX9BshcD5HJ08xoy9
4RZGs5XcCbHUleNyCcROolYSOHBqJUl7k3f8GN4McGx826pdubPBPQ9lZ0o5DZFi
QjMpBJupS5n5QIm4krbsavQSAjvOvzIjlgha4mWifPx5dzRsn43MncLPMIivRCV3
E3EO7LEOsbnVysMJdiHJVtMGWFLTbxxxf9UKKUFlcVJkKVr5vczvu8QhMRWqggzY
Gn1dK+kv7VaNjgs+B/RJYcUp+ENG32XAldyAm+mklxLTvxkZ7UCKwOjDOAdM+xEc
JwOuxX7p66Asa9XwVIfMqvobqcezubZk7pGIDhWBL3uBBuCN/JbKcijZhHXdnvaa
TfUi4duc/SPAuUzbfmVie6Go9DGMlPxKN5O/fA/f0cC6WEkI3LICsjyMX2CVpU5c
+n7l1mxX7/Ir6C0rttrsCw5pO/rbxgrntGakeOTV06N7ybDT8SzO3NM/C5sP7NM4
BqIgecjhGeUQIFb+VHrfshjKrwpOgUpfZ28mVAvuvO1XNmhg8/dxFXNjWbPya92f
dwjmHYNeATXQUOYtCRPqOUMXGkhBfAuE0TaIJntVDaAn9Nea+w6QJhV5ginZ1djI
tcBWKq/nnmHQ8r1q2Na5Stx3Yyd32asFXMcZLN8L3VtsjZr0XvakJviHJibAU+zg
GktJvqvIuRUQ5SEsPJ8d1iKsvSPsxYu16p/4f+3Oc0vnX44fHGAyJ2Q1wuR0xUTX
pfPNS/yb35beRvF7UavDTdnt35uqWAdTkCEG7sG7aqkcpzoL52BQXuoNeX7mMjV1
yIpNmvfK1zlW3jP4JqEff3akT0AkdTfWiCWZEGfZwYDDLOsU+URncm5NhrdVTfFG
K0zxivMt9PFHprtyJJpz/9leZ+Rw4lIzI8DqHXvsQ8ksVBoB2nqlvrcVGfkFWG/z
5rNXI5cXRRXsAv+xVRSLJvI82bgGVqCaI1h8iWxR5cS1CPrr5YZYttKzOizauoX7
Ru8spR8MNKM+n++dchWzLQH8GCUcBO4TWhwp0jQ9zc9OenDO/f/sLjVJqhh064uC
n44b+7D+kdJ8BGA6AdFXDQ9JMU9fSzC4ahZ3eEjAIbRLSLUT1sTohY6P397G2Q6L
Gb6vnFxsBVfRkKqty+CFSoFnl/62cOKPTZ26jezOb8g3nAq5vsA5kpgu0v9s6juQ
ta5mxaE0ydgZ/AAveGxubgJHfzEIFjLnogZu1/9eohNoqKi83yOHAVrlwq+6N+nD
CfugMH8Xbvfdn2NsgJQSgs7RUYdHpdWCTGixOwY4q5x1mm2YiuCwdakTUcK3h3jd
9stVKtbYU8qPooYs0NP3m6Q4Kd3Pv0RFZ1gNuYkUYItxv6qhKcNalDVYPzzybIs0
ZhPQklXZ4AJ3uzHzKptCCZpbWvr9kuWSFDaIIjyPcv0cbfuZ6dxi0/n6P53dwJW0
t+gCcoQBW/waeRiYgAgZ8uqRUcqpl/f60mUvq+OuqyjSstantxIFcBH5UHYGJps+
tT3GXxOBSFhVeMtCU4TcPkbxDSoCKDyc1urFz8P+kiShZuQIcTYc+ijMsPG9fZfW
9SERScNQWg/owyrwamiP29sUTC4IgEHimZV39t8AEMXFMzX5gl2VP8Mu9DvEaTDk
pH8+jIiK0kScouSQkOdSzs5PwiazC4Lr/aCS0UTG7oRNEICcNUmLG+N4/YfuTxt9
bTXhP0FGYKVwk5omJ6ynCPYsBDBTuT5Of0G1KCPYAb7d3j0GCFdkxgKvSsQfUfGg
+ii4MgUNwg0NJ3+eUoQrbr2OaHSdY53voElv7yWsq0U5BTOVzy1rIMod2SZIOeHl
Xps/M5gqVj9rm93ZY0R/X+QqkkOeVv8BOyBVkbATS5W1TxTbu+ywLvH2mJwM84Yt
RPAxvjLYbsKgdN1OXeElJxJqHq2Zv2w4TMFXSQardW9257YExFIPvV9m/lSzJGiO
+XSGhS/n25cGB7OoFanjhtDzsFb4rsFBU5v6CVdY1nxSXmBxqtEhLeK5WQvQfa7k
RIchpQaamgBTYCQhc4YtMT+xrItntJM9+mnuks6D3zptB/lI/CmLFRJjI93P+j6w
r7Q7evTuxol3++Ew8Q7rReNMkQn9R6oBc9Z5E1PDlJtypnE/wNV6sK7OF91lw7t1
Ky3KrVpzXKKfGzztFaQg3SdWaR+O3OWUv1ejtYiFNqbMEcMZEQTA4Url6cKvBFjG
zhNtYjfXQf8G7YAp0q0BFVWAe5DpLfu65h3cQTyRu3sLAG3Tvkjj8Tri+zKCFWcn
UqoIv4OQRxrYO0ZVNT/Ijpqf4WHP+KC/nNzYAtyUNx+Gn8rvgzGVfzUVvGmCRQVm
Hr/xV9+oskpt4oCpO6rbcm4otnNxSNOhkOPmIThegXWJbdfiuzIPnEz9wpqmEFpz
Hk7a+/eK83jblg34Cz4uZvGRxzPMEUXmoOazonOWOQLElendonaGPpTMZL1QgNlZ
fIXRzvxamja+tZrYyrZz5pfXC/jUXAYEhHchW+jOtnH1/ModazxpxpjrGivfCYJk
4rbLiQzkgzv+c1xpiEt+DFS7CLi3aOGwtdrxy869UP+2t7XwAeRPZyD0dge2B68Y
+Zhky+NtmRnrezcZ0pFmxJslfJPuxXFhmxVdqxJFbQ9WqK8lIQrBTPjoHsoj11JA
z9po0wnJJTgU98EUP+WELGZkTRyQUbDt+9w59qpXdchv9HV4udH2tAB3aQoU9x8a
D4pnRo+DJpaYSteEAxXxaxu4w528f4oLI/aRJynUlE9XoigGX2uM7tvpYdQ3cwOM
DWgOmiIIDLj0FnAMnaxFCfDZy0TzJfWREnsmROIkyOL8A/dPJTyUFrgwhenWqxeG
QQt8xZS9A/hcpA8rU2eSqChVYzJl0eTLb8uxkVrnikGCqU0TpfRvZrTZlIoBsYRl
l7xyDeajbTGh/WxIrQ2TXCI+oHo953VinZOCl2sigKcvj+elXPz5AVacgUL5efm9
QjsWCEUfTCVBkHJirNoq25wnrnuCb+1KqOOOlQakMZciH6tJyJOLaGMcCZ85lW3B
I+GD2Hk6D+MbAla/CTzazzRidzP3CzwycQNUsXPcmlkri+RGCkBqZgCMxLVIghOT
9+oqd06yzCSeznBgH/R7A31EtvcGHhlvfLoTHEYRXP6OIOoT3KTH1StUB/TELs2g
OqUzrmbqYxSDOrMlUHSyFzSyF3JzZw3vDgH9lOcBwAuYMHh2gvVEwqvcKEK1mr//
c0FCDBlE7MDWPA+pdiK6575XsLOmahpG0Ozg7lRFCbc7kD3FiEuWNA/VTceUPZSW
VID6wOD9rFvhNru74k+TG87JJsnzc80IhGyQVa1Jj6djn14NiTeANuKpxfZx3D2D
zPoiD5QqUSg4oU9YFQgMLu5LKHvSIq4m5lzQMqE+3indvC3YMCtF0+JZrMO/iocV
Oe3+fuvu2Yny4rmPuVhJuueSwE7iB8cnJxhsiZi2ejTjHa5Ltfs9ZlTklHWFBrBp
h8tAKf5Txc8TF7XWS52+VRjPnvUrcBd9VrJ0xILX2pSl6CTecOQZxzR0lymhUrQP
gy7x44FAiXiHRY3t0cJ4djUMqSVikJq+QUMQ/PeHjCyhorEUz74xt1bZFfbRVZ9V
xPDooYTtgbfqV/1P1Vc8q0Im/oTtiFsQ4Nl0L+iXhz181jkiSG3O9wduRC483xb2
ho4I6uNTuwABlIohRP5O7MGbNgd6vjoa6VqpsVnEjOn16pz9fS4uZ0laVgQFQyWb
WQKgtjwpi4ayObWMYIo0kI5mRVWu5bFBzIwcV6RgfPnWySd5WGYQoCtjx/KypU1z
g+cbK6niZuytxTWqzR4bTp5cVHznNff48ximF7ihvL/ZXuhtEEjno1HJnN1VCjy0
xv4EvnsIdi2gqdRwRQ7AyifuoXw/0bzYezCSG/AlJcNKGgc9x6Lbyoyapc/qGFdK
5Tat/4HFix/G16Xn2vI+9Wx25e9nfez4Z5+twugn6VlyGN1T+uG2dFfIuobGjZ0T
VOH8rpUpici5CB4y1CUUBQeJQ3WGV6fH3o4dJXiqYO71+wwnIo5+JBDNCt1vrKXV
hFQ7bfqKqIoqbVl8z7lWNthPggW0qASLVRVwA8dmMIUgQS5b9lLG/oTmNkVoiu4G
3nMJFQKfkbhWLbGhUl5cUoTDJywEjafQUx/Ue3KXUb4N/rspFmMfG+rIO3i3tBgL
xohqngW7hpTQ2+HyWBMo79h9meqZnS0Ugj3S74BE/tCeFChiT6Gn6skVisPph9x+
xUWo9HRuFFVqACSE07PjJgPL4WqZbUAokA7Xmkt0MOp6PQCpKjJKWbcBPd+Asvuf
KpGPeolTKk+sDXnppCTQwlmxE9gSIuYAdwdM8y/0G6qEebeKzIFy/b3tVXMHagU+
UZG09rwVviMl8bJUxRAt0abODeplrTTCKF/V0vOyHKTT4vYGvNTr2OZy5zfb+fup
YBua2+CEc4/UomAngSH0iUDxHVG7VXW1LtqOWOcdgelevyNtCw1YzDzcYsGRxvXF
nadQruGRh55RdSM8HkAGi+DnLKaSI2WOxMqI+DYDV99JmqtGCHpdt8TPuOOHLE19
WHrCqmONFLwK0oH2Ku4yPxXe5lkc3hFIgsggg5PmG89hfG6QP5+Td1AdQPn5UUsv
J5edscUNLXNSUtSH2xE/e1ZDYP7rwDtYFbM1o7Fx8uvmDQR3Z0J0GzFcMWwKllzw
1b46gtozucPQPPY71gFiiQCTi/lNEjCV+llc0bb1w6KZwPJvNy5tP/GodYsZfO3H
Dq0sfrOld+wvCrtwWHUYH/QOxe05ZoH1Ekl5bGD3AjrkkQoKiyarxHvKz2RkvYVC
o8MW+0e6wmK9+eu5LaZvjZtO/P8N4I1c2Txlk+iGUc8TU/DMSHe811/GMIlSJ232
QAhqojPM5w1/RTSa2pgv1pDbB0w4slrRj6bF+YT6a2rJtst0jq0j2sSNgE9XxZYM
zM3h8wTN1vZJp2thMwCqyc8Ag38NMQ22WWsQ6B7S0YVTeTkzcdxT4DSiUVeamVEj
r2YW7YS0aMr3kwDE9Z+jFr6JX5E4CvlLYyG8j37izDEHlzRv4qUGMDJnR16XWu1f
jVPQMEWMoceC3mrKuaMhfLPa3x0K0TktufAxfIFnkRjNDInyKzkI5X6bcPG7m8V7
lqT42ahQCpqvRUfaHShISRvqF2B2gIZ9dgZPXLiHMc+CjS89DS69V1QiVgXWni7z
/7hKyGt+h4oOX2fD3LpVle2yZbqDsJjJ3lfUeuXheIPoWwqyVjTEqjz49p+BFQ2I
qkZbskHY9J/cnZJSUSQADcoBEcFXt0BxlpivBKzjiQ62A4p7/lEwye5Xmp/KOSjM
BfCtjWbEZtHLA/HnOvOFAUnIe4xrdEceGr/qVkQQ41ZPb23rupHVeZfwnUT2XVPj
yJOpWdrNviY3ih9YT3JKXp3CNRieYkEjqfVzQ7Aed2XreP6nlpa+Jb6Xme7GAgry
NVJG+586u/EBy2UStNgfzNtJ648ITfMa+/Gu46XezDHZJ1tmdR8lrv2okHotUC6H
mCa7vnH+g76SrdYbEZkyTLvH0hR+BLdnDyWcKUD5ee3k5/Ohj3+WQKaIDbC/RB+5
OKff4kySuiKn01AX2NQV2srR9iFQBpXyMTYkUsLq1D+iBMUyT0SY+GFzAu7gSof6
xzznOIgvpZrfIu8jo6ZFNTS0RnGTWBtYU2QXKbrXCZ7zSlXnL4r7jEYjf7lSDfL1
IjcISk9kD74v8hbMj36d44J7M/s3EMjT0xGGPMgQw36Cx1GTNc2BBdQiD84PGHCe
QHOIJgRcX5hIrduBpqHl5vHYjMvvHfXcYh42qNbBeC9RnHo4wGV5l8VFXab6ojMK
h1OWOj8sPZ2CD4xgsLdY2lEtCN33iDRpxcGjl8GnzKqx2sSKxcAEShICdleWRxE2
fV2eWdkfncbXr6bOfZjMQA/GnMJMNnYm6/7cfPwYxPWf5Tb02hNZyD2wqnyC9tQc
Ll69XmnlAoWexPz71rBUiraj4LtE7aacj5DNpm29iefGUfSPswZzz6CHsGQhvj1R
o84LrkTgTDfNJ1SUjG5WRykhJ8O1luJwyrKRp/7+bxr4OWMjVNbhfsThwnT1vaYD
QS3hHmNapIdrMjWDv5/gLrlZ4YtY7uZnseZWPRaHyk7YJcjI31Kv6QIYiw3HXaHJ
W2Gba/ByS49HSCbkc9iBWOuDiZ8/RJh/SYMtfczANPAOTxk/KlQHa3zfBmXlPCWC
SGy9ZKfytt0avJtCy3tC5RuobsIin+y5w/i9MAupBJQlwWD3lMwepwKr21VA9VT2
Kg5oF1Qf49m4WqdToS2nXuG9mqIEeZ3oGXCHbeXFpTO5MZ1I+Kx6JeukSkqSEUuU
JeKH3tPPZu9Ea8bnWtkUrMW7jGQdqTZbmr+FcwE+M2H+BFjh4Q/IEMWLZEMwq1am
bfRiEh9N1Q27XjTotgjiBNKlkj3+uIvNysGX8oOAFfW95iFEb/OV3qvm3Ed3froP
2ozR1suRnV2HB5w3RixQZjDNZzkTs+uOZyxGZFAi3/N3EZwyZeMLtTBj0Ktw/Ks+
5Nh+MHncGCKw9yLIg7jUeCiXUcRcgLgjbT5n7+eutgNIRQqLgZDdRhMAWg+GqkPv
PlX6UaZ/53D1IcaxrTWgmimC/aXEcaC8y4fd0FX31whSsVyV+t1zm2vh0JYcX2Cq
IkEQoBeOc+xwqRVtlSN4k7WKk/SF2rAd/VrJ6UPtLGQXMK3wgRRfhMsur03zU+M3
iynnGDj2YnDX7wix8kmY5xeFgCOmzEa8lStedO3gKcctUwuVNaaG5e639tLQOHta
Cx+PguIxOMXB2RfPY+Y7L9DQpJRURiRq8YfbcjtgR7J9q4Q5dSe64ikhcVPEEKai
UvDE7veWjT5G1vYzFajX2l60+zk7cGyow/fswwnMTovZuCuguxBXAl8kxS9WxKPH
7E0K3mXa5IE7Eq01Y1JgNq4pb4R7Z84q0YY6W4rioDkpPh3+EgA1csDQ5UZFsrww
TgZyWngNLjrrExbt+snMepIxdcQ9o/5FTu+5clzOEtoHda+0rEH1oHh4AYPNfnCQ
fll9tUv8m7p9PMpzNI5Lth/LZPX55kkSVASz1n+/7c+2kuQ22aLPek+gdlsP/cPP
NUDC6abtaBlJQW2vuB1cIVqACXGhanCIr3Ta19vsEFkN20zY7HhydQbnfxu4DCOJ
GIuzF3GiAbMiiHvf8PLMkvf9/7mXQZI1zYqQnu5jf5KfolM7r6I+7dHCe7t6Mz+U
HRkx8jNP9rqpG5xGONa+vA3x/c2WOc2FM0UzZwmZ8oYvL0vdU27LmkXh3/rs6Tu1
Fv0l3ODxTJeta+HKciSS7tvjbIWiZ54h2TvzMIHys4oUvtm5QHzgQP/GAkNWMrKQ
srywNh7eimV+jNpm8y/Rkz39NjtUYq9hOVzQZND9cRLwuFB8yrUtEQbGUltJDjTR
7IBJOf/hNV3Jxfwelzj4bSLR0E18ryO5r0MVt5Df0zr0nUibKUepf2/gFfEcKB1J
cx711cj8QRn3n7+LNEO/wFRBmkEFc8lGSgKQ+5k+Y9fTEQYU8fD4znJIlQaaxVc6
V2wP+I7gncVcmC/C7Vysgsg3IZw63jKjSuzlQt9LbUInzrQqeuXitkl+KJ+ZFx+M
9pVdX85K3W64kUguLub+P6xboVaUmqlJ2T0LnzboZ7QIng0LvFqdXpp13fyoEXD1
Uo11usmzNEl3V3Y7v58VOvozCs5cibm2DxjHk8oWO6DLc0v6ESFq0wuHlxuu/bJl
HjZ+bzCJsCzOMhjgrTx1ZCnH34lBw+8xw3zv3u52XCMiLNQ5eYwLuE8Nnfc3NpN3
jh0juRXex1R4aeHskWs0Vm6z1opbraJxR3g7G6OVyhLT4cgjRL28IfLZiTomt08m
u3HU3z8YBApipSPmT0DbVHoxmLIzCgkpv88N3GgJDdiQY+OSXDAeJqHAvPBI2gjw
67sJqLcpO9oAONEKhlLypKUB9hcK8+2/+OuRDwppiPoFc9BcpAMVJX8faD9EikP/
Di2VL5NfIMyMZO+/SzyyMOn5YKlkxwO3yXKQzROcA7OGHjKdui6TLX3TQM4xuMAK
rC6gCr7m2E2kKIBvfBaZiqP9hgIWVumDleMuW/hOQPr4b4QrMS1aDmoAq70TW2fH
pBhorFr4ongM9Lw9u8m2US/WsurijqLAwTcXT77INKPZlRjXK23qpf4B0queJZZV
VORMWUzOgca95z+w1MLKZ8Vx4y/afYLNG/D6FevvlT+T3Vtzxj7wkWqCGcOyrBY0
idE1AY16B51kDT7L5Yh/pLfrD8EzHXqmh/+V1VrfTbUbLFb9U/E7Tb/qUaAgAEKc
CwtGnOi+nk6nq6AieSBc/XUNtQoRcz3KnW2OOQrwRotIoXzvknxiwXUfafD5kdZp
iVWntVGlUpUFiricXFM3yKIjXt4VmZ6ILFu4ecrvK4esIySK7TfRQL5JIbctxohE
yhAUcXGCTb6OeO7F/153Um/d7y36JH779pa6X/5QqudzBfEYOkDmVheg2PW+52MC
9PrdEU1bSIWx/X4AdaD4evLMS9QevwWMUFqLzubtDf2dapOLvZmhL1D2aTstbqdk
AbnJ62eDTfM8R+Zyn/I0AVwwsNvN7ZniVp8MhcAI77JStnyEx7TOLueqGcf85cEz
ja/mv6S4uCuuVMc5F8KBMCPhNYVlI8E4WmeHywEYUHn/o2BRazYr247lquW5t3KJ
F4E6Qbce6az7akwiNzSILXcEoMnRJwNe1t1g96cygT6kAULWPvCshbTHkk14qljb
zeyn1YzNP+6Y/nRcuoE+hMLhQ6AfEC3Ruo30+9wHGa11eh96PneoZA9ujzM+JqwV
xWY59ZPeQm1JpspcDrRhCgGas7GSy+elERqQuM1OcCONEQNGRV0NE6S7AdAXjgvc
rxAZr1nEDUqIeUaj3XLeVjhsXZAFxi9FVvjTRT/AdOpAPxt5pTLWOB+elKg9dus6
XcdMCXwKdfdEwqZKhOKuKpm9UshkzPZbQdPxFWdnrYpyTpVnlLppgeTFefARjEQy
UD6YubAzUi8AbaiqnIlW1oz1/WAnE2dvFLSLpQ/Al3ojbNkAE56fNDdhdqe0J3TQ
V7wBxXO7PtBm5aWSX9MF3HZoLaZDBsrc1BspwU01T0QDMIs235hSGUF1vFeHt3Li
VC0uVQHMCrVbRm4PuzbQXG2ezUUbOu2kZxG/pmq0MHTDhTfgs4JvzAP/X1eMGSW1
luAfAFFxGsy4UF5vIvXT05Y038gxi7kFtrOQauS28iS0SFVC5UP5PyyYIIRkWrUJ
nJHNRN4wX/eRf5zfluVQP2LPyHlWcn1WnJX+KW/AHtq5h5eFlGlvBws28zZPmkTW
eVw25LVJKe6lILEqClYIEX5KHaysEb1f6GZvyR+hJ7OAqNJ+Hc952Y4jMWNcs/Ry
ziH0Q/4mEkBWu8ihl4pWwOZhyaKzzx1jfOvYUQYdUV0Qupjgt/EJzfXvI7G1miOm
STdTHDmUSX8Zku16Zjk5T8HolMgUwVKi89PeU6YrvB8labL4u+TGDNvsZt5A6nzG
iRbNMJUWb41qZlGbvl2lU4xIhKHwNgjy/16TP7EOhmZE5y+KXdC0ZJ3D0mFjp9oc
PlgaF1vY8zf/3QeGMyXW5XBKgVtOp+58tgOXB98yvLcay+GWIg9ePOgyCM3ehPeO
xIjWl2SU7mqf11AnSuevrx7ufkCXAfvjWa5iBXGx0E2l5Kgaa1FZpiILq5mIkqnN
bhSAQ+LM/5aEcqHt3nLiPyj1VtKcuHKFeKegPE9CLyVcEwtaTzWYzTTAieEhGerM
JjUWqMMX9+JqUK3bIUjfP5fNkVKEiehBeh536DL+B7hIKWYr4ABvyLouygK40HZP
wKaANUoFAgF4sekTP7xdQl4pYOU4U5FjRG7D55e+a+0I8tly+0EBKqXuExypsL5k
lKcoLsSd0rJjtdIm5yRI4VncJvjHwF6maYTJA0LzwUTIiOnYSxjqC6StETmkYJc0
bDC3OzYn93Qvz2+6upl/o2PcnGN7V8yk7UzBx99XQrssWZXsxNsQGFMWNukbp3Yr
eiIewhBm8Qmql2+KVBconbHyE/bo44rfgJj1N0BP94fI019hvNfQ7USmYHPMmgZ6
J/mw2/U83ke3ptI76OGCR1dvzv9g066AssHPyBz8GIJiv64wNJjTJs54ho03f6rK
3fQccePS//6S+zR7osmbsdImnz2nzJbJFhdRZNGwKNqbfdFE8E4r8/o7KcRpqoc7
l0TlikL7GnHdzNsy57SEtTXYq21GiVeeK6DIMHmftD9IWthrblub3QmHCDvWOqYA
2d7dk8kR7wYcYSLqBnBEDv7MOuBJ084Cppp/fYIaWmS4hQOOvfp6Lp0oUOL3GL8h
4hJufL68XUsfzYOG+wkiH/njxTa/OK2LQvNT+0kVJDhlvMXTANks6j4Lbm9p0Lav
rzHSQudpJ4GYU2ZTsC9oNHUF5kItV78gDLlgEIFdPb7J2RJk39nZk4SXWIAtP5kw
NEx2zqy7fecKgU4PtTpDTkFWEPJzH27uJnx1TpuofpPqY+fkqXm3yVlYLnIxRqua
k9MgLPD3eLqMRyTOLGWlupa710RHaJpHtgq8QeiMaxHL2y+sfCMzTUAFDEFxEn+I
PVlut96UKRlO0a3wgSTW0/Wj77sJH7weSewPb+YKZcQP1lW9G/Z9Jb1RU2MFSJ4S
Im7LI4qE5sRyDmMGFi907Y3TBsGCtmQvwnqV8gykYNWryvieoIZnAePcuqoGxxpP
VQPb5tygE2VVOleKQLKnU8h7ofcxs7jpTzTiI36g3yd8mqQLeRETRT5NosCbYNpW
wwuSuAknkoYtU5u0QXhoZ2meIY/cpERTa3OJcz+sGMXoWgUQFhGVPXxYwVhYij4o
o96UvGHtFzc04W4k5BoMhZXRCCdawDuFmTTIPlVghRmGSp6IbOPTPWgi2Qm0MREi
ms8Ij4cIBWp7jX+HVgIZwZZctCT3p9LxKyo3S+Ji7GrZV+CBSqQR44DdS6EWx9eO
TFos3cGzi0wYEpVcRlTYCyBisUeJkDhQKieSQT25W8lG9N8xVEEN+ICeSt4UiG2Z
6g2MY1U2fyIKdIzSUE7bPCen7HH50DDrnnJWulI22JT29uL/dcXAPCabDj9BfZ0h
ct5FcTAY0iIctEuRx+OWhcKEXU50SaYXJDWTyD2+B0dxtkbGPpzdpFjQomiPkKaH
xk0364sIGE4HcSTP+WEIcGgFsMCdz66y7cpxuJwvehDAfshlCKom/9lKdzm27T3F
/n3621kjrBgZyyWE49R5XZ8/Uv7ES5MqfZ8bMaRz6CWmql1qNBjO8J4zCgMkPWPO
/lpmQcsUeCaA+ugSzGKAiaF0a0jWsTMWAcR3B3/jS42AsG8StuQvfPkWAWo7qU8N
q1HW+OmHYc2Sn7ECiH8Bo3fKnVv3yeM1TLSTF2BMB49LJgl4g354Dy4x2uIw2Np6
wCwSN6wAawMrFjKWz73aVOHVRzZkMluT5yq/lA1ErhB588T0eE8uTTN9LxvVyvK3
o0T3tjp47l6NGvwijcHoXm7DEIznx48fXTcGRzerIsd4wcLSeRefG6v36hHnMSpl
wWhHWfu5CuyvGsPxyVf5Ld8N2IDy9rt2C1/5iNltbvTxiNOPxlcUQKf+o5Owl3Qq
OUwQJU0vknekzefdKQ5qiMgw4rHzUu3oAjtXE9gXKILT8zmpsl7dj1h8aX0HQXp1
a0f6xMcXrvOqSqrSnl0nmSQVggqIz6n69UUTRh6IOnAIjlUWKACaiGJLIhYEozqg
6fMZtqfMERqlNbWfdakvA7++rjRIGPWi/adYhz/rmLnDogxhjw+qPC4FatlU9SGb
WJG0pHKnc6IGIOmjzqFB0VtAmcN4wMP/HYjBFr3sZENVUv7e68hYeQ6BMn94OT+a
K8OSJ7cJM8XNXhWKD523mOifwsVyTmu46QTiGzSK23hA8Ay/v+G3STFFfgpQxDjD
Bb9rKHaSmM5RL/yjC6lxwh/KEnU4BcZX2B1N4VHWyGdBiriE0oUBHzMKWK/VmMAk
1jQo2ekJGPu0A2kRkMjg+XW/dXD2s8qOvscRoatquLkqoXTAXskd4l/Cj+8onpge
Xg7+YI7s61IMHVmVA7dmnV5TbX9vxtglucv1S302jaCJq0IhHpz84X0rfRJVw6Az
FlXGwnfuUA3iYF3rYgyZPUPDPAGipmvgl8zVO1GgjJ1u8PkhqEsxDRWH7fOM6fla
`protect end_protected
