`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
O0D3XC+qDF5c4qlm77cnwf9VgJAzi/sfsul/57E2jIThpx/aU2u+4cqeki9mQUdP
SqfyrRTpzL5BHnby8fy5wqy8VvNdxBuHAPmnPOEVIclY36XeJWIiuYDPjnBDuGBw
dBSrynaYdPNZ2d5GFcwbZ1tk6sDgwquAWF9AM+Pln4eTm84VCrPa2Am4lJeBIps6
W8HivOr3E3AFhNQHZzP2auQbQo3K+96EHHBNMUvSEW3wPeADb19CLAw3LL9sUpJn
mfuxEm7tCKdp349eQTilN1O3jPK5m247VDv7jPlb+tc+AYFJxptbYMOdQw8E9Y2J
//zWyfGfogsIuvyT0yjO9w==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
HRXN3GhdsTp3rawRGGCZuLvirgsmm2+emHAGYv8mez3h7vbbC4F6C/O9qQZcQMVz
o5arEPzFzkkPN3rNbHVpSBsLKZz7bVeq+jUE/ZBMYnjQcXl3DRpsl09p4NXyvEKD
8K0rDOcG/UVXLaVoWqHQYiUrw7oFE3ZdRxVt82HWtGw=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5712 )
`protect data_block
jayrEIvQJuRONoy9pXULEf7hqFrOhbGCAu+EhNR29iLYNxH/LBAuRMZUg1DG2w2T
soh1Z/wfO8RWQXE59d92os7tvAAmh2T/Q0FyYmU5EeNKk8r8Nc4oLQWS/m/LAf/5
qkLIE82NxlfYr9WdQPYtw8EfTMyWPWQbMl8REmyajf5n4CALn1/x5YUfOLLV1Kvh
HjvCKmXd+vz9uV4Jr1t+V3NUM9nomVhb0gV/nn86BiLM29HwUH31uoDG5py18CnY
yZT/gqVG8UcJtpspTfh17tLB90PwJIRT8KS1JeXijPD6tyehVUZsWy7drrQSEHtk
chfq4VID/L8QffblX6xcu9VDfaTbTPAc1lquverkJe2aeVRq+WudCyn5+ibbNiwS
NkOtKtt4Vht7JkFU0yWd3ALibD3oiY+G5JChUgvt64Ur6HGhw2IZHPH8dkplB/BO
1OBnEalmpprpnWmlqJjxwlUrs0V83Rkx/xt/Y8DggrQG7aBhRnx2GMHfnKVqiFfe
l8ndo9q6TwRwth9SBA96XXl+Y0zqJ6wj5c10xJnmHDtHQAmatCMa3ozknjFPVewp
6RK/B84/Z5R5aRcnu+ikS/O9a7Tjksn+2AMn+jbofie0p7iVdcADCLc00/Ccf5Ru
JLgHCtuhPK8uDGbY/lqsEvYwwrxVPfeJuj6dlMf8RcdcyoqBpTTVLn7eOo+ZoEw4
k+wXLvtCP2lr0gas+gCp+Le/XWLuR6PLcYHOI8sDNhhkq50Ahe8bNQtqUoxYNHYj
6A150q7i+PGEYJZx4zYnCruZTFV9+QV68MMSulKEKwbu4/c1UaO7dqPDKHKbdikH
r6bBUODOxnZnGg45eMHbZJKYYSrZZxqb9wM8FjqNWuqSyj3xdyDapR0sa22kBWW2
W11eh6YVKAyb6kfCVx4BvOA0QwZp5UvXuIxGGXZwPT4e5dZEAfqsfo6QQvk28LZZ
pvTpyj6OVCjIxpfmy4SlkB9yHvJJHx8Z0ciqHy+ku6dBv7JPF78o0Dq4Ww8U14lq
NAQTImPoAVOphfl72Kuma4QXJitYS9Q1yoPkq+I5rhXg1njvFmmeG/JtcnLwz4cG
06MI+l9bq3tSNVytkfvTygRGaqhqOIIDKQhcUhGqUTOibfMOcA0VHtb6BuLtRQnv
ILu62QxGtMDxqogYYkBhscOR5EHcLI4PtcZE/zRCFzQBMqaVauP01PY/H0Kxcck9
gRqD1q1T2mHOmp7NSSu0ZmtX89uyPEf1nRS6nOINTyL8Q49JjuEtwiNuPQxXRUyt
dXRXOZsP2XCfEtCwd4GOhjJo0tvr/noBjwU3FEFxuT+7Run9KQrVSbqU+Em7wj79
nMNmXvDmLLiciZnsEyisO26zanFdreHknp5Vsv3GIwpMMI7n97LnIhh7gq7ukIKT
yUjrtHCwcW6hc5AhSnVSwxaGMKS6k697t1lTwu78S3RhiVo/xC31ycZqVKOUCrgW
i9dWcu434y9ojMtgkhnlxGMontjINivzbU+1BozmjBlJvJ4SjBxqotQUz10DFag6
QsbNSrc6eEFhVhXc1XDvszW1dryuxYGgkDS9pf9MixRFCEvwRElekNhdCoVwpV8u
B1jZ0aOeejhugPtYmdSDyxEgjZhOxMHaKdFpBf82jtlap4RlXargBxGe5cAuUSRN
buHtljUZ5gGpSRScGKjnZ2pwgUVTIDfvOPTyN+CzdJ6pnAVUM0LVRk7u3e8ld8am
QdFIOaMJIDwYvXvgWvW+NbjNFi6mgDAKZ9aLmvEjy/EXZNW3scwViZ5JSNq4pGZo
hBmsG205wO1qv4eEb+ZxYSof0tbNt3GbxEVR4vB3gHSehfESJAojhFOr4RSeMui4
ILcY7q8wL/N4qo8SJ2lp2uO8gNMiwaL0L3DwqYwJo0HYF3EgQjXTBpgUQ5MNJ5Wp
G9ZxX/GLMYroY2m0el2ECYnZJB4/rZuBYG6qfWpYhx5oIwdoGyongORvzAHM4Ynq
2Pun16Hi1DigalVyUOYtfJ4uDRpRuhhEu/CO4LRcCU1+0Gr6u4Pt0Qd2pR7V/IZF
mOkAtyUDl2xRDd6m6kcuCL05+mYtxIRwRAMyc1BOgoUUgYFX5mYxFlUBiijmqu6i
mzUvNOKlOqhWPteqKePUbDAe5Da4w9a4Qfdy6p1F4fBPakgaa8eIpTFHhi1C6sZk
hr/0R5nd1ZpHrohkQ/CEDsTBMJsNLPPrCcAxUJStjwXRBvA8mBIpC6lSyBWqjnaI
KCXCz58QAXbt7rIVIo2oFzOc3m0aQB5JkC0YQPIzzYVQMeekAiI51OFpzXEYLuUJ
CLa+IvNUVPPu/tmm5t4+du9M97kRP9oSerFtSVnyNo69UzJ5WdAxOd5ysZUqStAS
P4s0LFMKyUk5zjXHxk+DM7z508+37suLo3w5gl5eg5BziknQ7dy/dkYz6hVxdeXh
wsvtzYXLfCHmS2thk8jetva+ZxY5BTm7R+Ra6ZYuXuKj4IjPrMIp2ndXmT2BPT5C
zLVqxlud7i9DNy3XvaFeUk7i1+rDbtQXQmyTTAgTesb//VNySy/LoDKpY07Jw8ZA
6aENK9dWcMHegqBDRAiI34gFEHXRiBqQL7JFbug58a3yaT9W82el3XHFijzmPWKC
OXUrsnVcNjNlRHe3w+Y3lTT6hf4iWhSh5BCj2rHcENxQ3JdRPa7bDMK/4txmeFoJ
mkPHzzObfL+ETMYhFm11jd7vmx9e7g6P4UaenP5YQZRuN/IYH1ZVER82dmnb1ra7
DN9Z0OqqOzTcG+J1YQGtfvXs8W2jyKaBTRQgHyPrGYISljn2scjhmdnbge9b6VA4
jm48Dh68z7sZBKKf18SKYvJIwOS/YFIG/ldMipIaKxFFqohdjveQ5hN8hpcqQI+O
Q3tDicd/J2wGFD53QzHjpPX6YqFuz4eXjklc0kqTLBOZTd8hC6VKGu3QNOnZJz2g
KvIYhDI+ara4NoTGAGiN5KWgAVEz+jtm5V3PQv2lSupEM74tlG/vMvr/tyCRBU89
fQD2jRkT1shXTYGETzcje9SD/VYn2LPSJ8O5PAGeWoraFbiqE7dBVJDInC4tvS5V
A/iPbT1wUxJrEYu2fYSq3XxgeWXvmHft+1XyGG7IZdq2sj8sUsp4YRnqN8pYPU50
DyvVN5hZ7yExBwg/t2zWPus1C5TrFwouR0kJKp3NwyyBIfwnpmJFuolS5sO25WOA
fM35nJFRb+VqBeckwSZ/1BxvDXEWbsHkZyBq9J/z/5CrVCtPg6u8UKLn/vJg8vjo
p+jGLKaLzSA+e++iPOVBErZ3wCwZBHj2E0K7jWHGAxooMVdxsWGfP3x2p8ixciQt
pO+6LeEPkBxLPF9ejJnwt2Rd19Rhea9zYwfVqsk9IYozVJKi18G4C457hkz8htEQ
Dm6in9bnfKiEb1Gjd4WBIgKZ2ap7v4UZS4ZMdsPH+TmtP0jZ5F9+5hjhNdnJ6/tI
oSjXUKXVNw6en5TSxWFhcwxUOfWb/71uWsxmhNlxJhI3xHW+0DD3w5ZXtGZFbuWi
4Jpr3MFYuLkSKA6UbtA+rFx1aLTOm9H+NlIiQpR8Mn2OPtvfN0g96NZX16KGGzCW
fq0/OFphOIP1gEqQ1yORGum0/E1Y9Jr1JpUv71ghQDJpFYwETplImdfsNiVmC+L/
uSxsSNOTxFJfk9sYQJ4Jm3dITYZU3CILwxIvp44U6UnzlK9aFyj/iZHxfRuaB7ip
IiEBE3nVvtjBuWqQ6kJuNz5pTlCdG+gDyU8PwFHf/t8OucW1Ki4QCoZqd7cN18q/
r/qqjd3p8xMrdDKE54ErO9esn0HhrSs+ULPmz8jfA4WmnRDZ4DqhgwIYord8CWEW
ub5CCLzNQleBgnf7hDIYTd/cQcOq08tG2sAK213FQLWBTQ0PxhzznO6h2evZl+ei
hCICNupfHv/Lm5XlUDluc+HsKyXfzN0weJn3ppPaGK4ieTCm1yYN4z2ysbLf+q3P
wlnVLoDpiudv9Yx1E4UgbRMv02+XmWD68TNB5tgARNRZ8jA7tBNdAwVI3ITGWaow
pfWs4kkFoq6TbLZNPqSfmNlutfYfHTC436gV/Jvg/zB7dbsdBUUSjn+eFwwwvWG3
yVq+PFB8KuEWP87W00bhU6MPWbKZX3Xh+b75zgB1VE6siAJZNJSDL7NuDNRcZZTd
S1OAOmMQm0CftBLNoovquUIDFgjxXgMPqDoN5CA8d/IkCPKfI8Dgg7SZMUUV2AQE
0PFQbfOL5ZWOXPEKgc9uqr7h1B+IsyNZJFF0tFaq/xQBo/sm6Z2UlMQLg+UR8s6f
9VszVeIyvV48oL1lMyj5LcEouVIEPWdhZjVFk8YEQQUSzQc8N4yTWoNNyxj3WAXp
054lUJZHI4vOx4R+TT/mYQhBp8vzxnzpweI+/8N8AzyREuR/iMAhMrLE7qDtSZfF
X0m0LzN/6N929AKWhM2hzcRhFYN3Sw7jOppxX9dFkrcPwi2COnR+8GVVDlV3T2Nj
jheua0s+uKvhmbmp2Nz7qxgAr+lhpP3RbGI7fQEmJOBcRv6seA1KHSK92cu2vtR/
tkB2A8KlzYxhbQGutVd3BhmA28tGyoR+05DYQr76C9w5zkLpUEx1HkWVKL72sen3
IjLhKLA7+vt2gXgAts18t5gdAe9VZZUW9OStDImc8d/cqXb3IEBfqfc2c5eLKhPZ
Ojj4Mj+aNBml0qBJsVCafg0UNSazNusohOYfU6X3jpFt1Y4exDTN7EQWP6pQJdNp
vryPtKYuFz9QAxlb4lH58t86qFWFh7YJbriCc+UEntaoGHT7hM2JqYhJ1z4q68ij
99Y44FFQ4WOK8UZj0hNoXp2eVbHPUHF3JFjFbSQQHHM45/GNyIOFT5kFyUn6HBHz
Sbp5EWdFGu1mUcdXeCmJu/19XYjjPDYuhmm8ikc2dPRzYyCSlOQ3P4TaAmQaC/NL
uzrqt0qKuwaIFRKwvHbcffWqM+NMdpOspn60g+9djBF/WLCftXtMjnrvrJHFmC8A
yqw+4xItCTDchf2iIbbcfUYhB49R2MbSyecwVrD79P59lkJ/904un/mQXcAGTRgr
Ut3MwC2C1uguA7Vypxz24NVXRQRLUQZiX7c71mA6+bt9L+e0yzIaSKC1ShMeRHDD
zFm3/QUS6m19Pn2IsOPFKDZF6FYOpqP6HFFo4BMWx/30Oce0wXdYiSb5xO9l/hId
26lCRtsp9HE9CHKCey2t7BD+p76pW5kycHNlFuIxb7KTsCsUrtxTREfDIp2lhKa9
Y62nytW3pKbRh25Am9u8LSLIom1ASELusfdm/WdDNl3kKlAU97+bWx5+hxZ93pQ3
A9fqV6XgRv87ge+trKqNnJZTJrSaOIF/y13QamJTcFbQlboEHV8jljVoMmlbMFKG
fDv3E0a4IcmkWhTm1UnndNX6d9iU4oJVoiPyBAw62rn/y5So2o/3apAGfWH74Ont
KB6hEE2X9ZquEp20kx50gvasJmH27RJYSHMYNastWjRypgYzPhriFzub57XNiuBu
DltVI0/yhiaCnehP+PdVGVTCM3mGsPhI+xBYNh8nfmhh8CayvC4a+vYmwb3wZgM/
Rf0oL/+IaWYYm6n9SKDhGy1QkDD3MwzP1LpE6bItcBNPQxm3nnq8/Kg41N39Zhbv
ws2ydHLMZK6vXfUw2ZBy+8QaB4OWAQ4hbvJTrIEo+H3rXgDSoSy7zQC8j2Ye+fqX
6LZtXZy3kXjmSLmM4QwUB6+bnMIjdLl13eK81Wfj3OW7Ajp5KmnC+wtoIkaDSp30
wHBFMY+9apjfiXJPwgA8sFILdyTG/L4ly8HaI7hTzxhltI6Uggq2Rnvdkb+1x0GT
6Bo9ONsi2s7FUZyVfrOTnZl0tLm3qRZFSbMJX25Y2KWrTltmFyozx6YicOAXfDhw
Pt8sn04wAIlXHApweIUlCOdFjZ4phYzTuSdafUw1wtHd2feO2D++Q9sbeYOAlRjP
CQlQeLilpGbygtaAQghuGfXUb9z6avkncohBby4k1QcsLFTtgencs/OqT4YbaVsM
j5phN39Mjl2J2PS0GexYYj8KQtjrk8nq4Nrbnw75QzMuXD+H4DF1sg2YAqsmwg33
Si1/2evCFtyRThmaoLCPQeplurz9UkaZx6svo+gpxZNW3nDtNK/+qwZFZHIz4cuf
PlKzSyGQVoI8yKV+yw/L7zSbgdMSNmPvHtArQrQTolb5nSUe0sIN9HMkQER0YQ6y
GvvuMSu0aDgLBDV/l8brtGUaNTosbcmNqcZOCh35EXR1NKAAF+nJPyan0R6jSZth
kusT0+EbXGCfVgU9sXO5uYdBRQRhmzAtMBVog8e96NC53S/Y9rm/rBV30EKqq0DF
f1J3vrZr1NO2F9/RblQf2LEGcPYZYq2sPahs32gp7daGvNyEeOGO6z+RpqB6ykHA
21CuE39rMNZX6NHxmgXsoGVqO850V4x6hE/mtDF8qKgZ9EqH/cnnGTB21nNbg1y1
tVAf061zKVmTlucBlS2gN5urb8p+AxCDw3EIvdiT75ep1O+27ASHEAQENy8JKx4d
du1tycG9jTt5o/9mHOnv5n7+9tx5WgTpR3nxhYa/SJaGPVYQ9BfNF9cD2nzEwgjM
l47btA+Hzwp0NX6hXrHtRsGMLOzaJaQyo3W6bVQarBpQ8d6vQHksCYm/kowlcVjY
YbngTjE9AJLw5OKXRs/TrmgZD0H23Wv3z5oY1h3LZxmoBNbaDSGOjdHonWuKNgm4
oYY0ELeYFEn+l2mmoqtyce0f0PqchuKtzbnNKcsfPFhfu3tx+jhQ72TJbjfr7NkQ
5zPuH3Zs7Oz+DR/xCbYWU07RpWq3JJ6xsUYY05tgKnWCbnJZaK6mZ1lee70T6lcG
D/41ysGo0aMg+tAgFNJEEQOOlUAdESsQ+Y86GmMQ1PvYugZPA2e5eoGoqnDjPHa5
7LsfPMLtC3yH8q7MvsHxtIaH9KULe4FO0nXgxRMFavCQSN+xmaDWPFmhJK0QV/qw
ktmEoZ7FqCU2SE9fy/MLqUPv4jPX96zbK6T5BBCqSNGXpZ5b6JA9jAZR7mNWjysy
Jpk/LT8vdmKPPSiyG5UYF+CTDU5J/fp7t7TSEunNcAJTa4ti9kxVJUrqukbPTNY2
4FjV9h7bc2QQztI7JGasCe2dHwddGlHxs5vSDI2iNJJZjc0WpUDbBp8wM+zLB5vX
aPNyoGA65Fch7+UWVrXKfsidRSWBd6lyk5sZmn4IURj8tFwozFog7FkjC+XomNNu
WS4kviMdzXDM+L86RuxDPs2TlAaYVrjpoLWKivmwKpVKRZlckecVrNW1WO/PKxY4
01JXdqhwqH+nSZE3l/DaWJtbuIZ2hCSEB2APiuxDD7gWowu55CbGWFzcyWNEZyhc
OHyPa4y9G72zvrbRHW2cQKRpWFsQ8osIhrOrrX6p3+TVqnvPOKuLcT2r7JgtfyKX
GzwuhYznYvIqHaKWXXFkYUq52goKRrzw88ux4LLipvYZ4CHk+fzefl2pY8De/mbB
EQ7SNylKbco558zHuo3bveujEVDX8BrFe+zltoSmiTkjlphWl6xdj4yX5R2ByFdF
WFhaifN41QkCmkkQEfrqXfc6p9tgtQM7uLYWp1CeS8dnRvgwcvVjsP+okhQtPt8h
`protect end_protected
