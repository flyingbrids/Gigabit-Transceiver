`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
o/k0lhxw21H+CtjYXqk0GDS/L8YvggaT+8XBCzXXgWoS9MfFFP503+13qGkReoyG
510xsgigqahRKUm566ssgcD6ehyCmZU/Qwm2SBAGR2FYQTJweHYFVlfE9QIp4zMz
1RSm3whKABTc+4PTOXiD45qo0lgG7AXO/JIZPCIivn0qusgxmFsUaNl2KgyV75Zd
d+4RJMPYVz6o7/u0VXuFNlmDfrO15ytWFvKVjkeaIjEjkZoPvHGlJAye0kLmx4Ap
emdQTBeE5+YFFQFHU3UlpxfT89+wVXUw7+5yCgPFHQMdqw5CcKyoYyGqqp1GQ9UC
PsV8emmPr3LoRLjgpMSqGw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
UYWNVKZqak9FlyI0HPunv6teIbCbm3Gt6mkGQ6tQHW80aj7iloM0Gf5uU9h5APGE
SE6xfbsQJIQ4+H4G1FPjn577Z0bjcz7GO4DZRzK+qONHS763qunrMdnXZMIh+6Tp
QOyVrN7sVvOiEDvIGx7aIPvmfz3OoLUFDJTqFql09As=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14080 )
`protect data_block
zKn+B4lfd1KAy2NJZdOjlA4VyZ0w7U6FRB3AW7nGybvQYK3gYuaCKmGrxTPNdiV6
H5za6IkEmmAcELyasXX5WuMPSy+BavOCWi20vDREyaCfY7YOsUMtuo+yMTRVr4o6
MhLxct31O40ZR3tJV2TxuxsawdMC3C5ilTU5ZITQivWdZON7tSf8niN0mMlWIB4K
hLyOyY4+mhWJXT095jZ5hTsraNudJkoExbNAeC4hE7kvRWixJe/myXLPkK1adMuJ
rAd4lIjGAUPfUvFYNdXzL6KKTDSofvEOXz3faSFWPbFPOZZx+7JaMbPsoiP6ijuu
rcV6wUZDV44rh4yN/TMVUyKQsbtrnZS7v+lyITGtVj7GueF/3XfIRK3E+dmC7sWs
B2pPHK6dRaxFRUVvSVvZGs9flYP5vZ4TKjTE/oe/R+AhxlJ598+Iw2fBmkAW5wWU
2JN4q/ED3kAo9qEns59f4ylL729u0B+2l0r+iGBnm+GMhYRhqpD3ynIkcGUwOTS9
kar+0umzrhrwXq2yr8uGWkZ9B5Osfqvsc7VYM7uBH7pO1LzHPOPdIvcTq0skmbPf
/Au2j8/ifDhyG5rqm8Na41Fuhc4zeoBYDF1SeWL2aW8dtyw4CPVRADCIjyxw8lbx
f30HPLBZ5nsJ15WrNiQpEvCZFY8sQQZJU4mAgZe1JHBn96F84hYusBL5Yss0737A
V8tuHQvnIJkWYbqdbNgNu4FT2iP8J1FnRluWLUjZvsE4TdEnJFTR0JTjD5XsqFet
OTJ9pcYd3BtY9fAmac/DOZstlCFS46YrIAmNve5meDJcygDSjraS4YxhTSsPbcl4
upHrwJgEWLCf1ijggn8az4fTYrAkeOLCJh6lJkpBdRUfwSsVmXiBIE08ok2M/CUn
XBR8LYlb3FqG/30AYCCq77ZQq7wbG8pDHx1MGM+JUYC998ihJudecXMWl9x0BpO7
RO1C8si6kwZcQIb7RNigHaRyn2Sme6PviSPWYsgnEgzgBpF1w5nCdDQu5FglwJiL
30Pr73XWmIZyuOGaDAzhqqr3c2uC6gBRGXouMMIrBZ4be2dE20Ob2gvu9msIZ93E
PQeJQMnPBtxd1PWZakqbccVguXU4ZzC3+ifio8JeF01PX+RFJH0eTo4kHvwzD0pw
9syZ4F+FUzBIU2LUYB4NBX7Cfd/m5UnHFZtqWZwZDzPVTwW5FvZ/2sFUfFzrVuJr
aDsAx3YRh9cxX/MsdrfQinEPzhso6yxBfM8GNJ/MMwnlFzg+ykUKA0/b2KOq25jn
jHIro8WZJs9KqQdvp8BW/NfxIcqN3sB3iBHBDXn0Ykvj+V4NY+23iAuCKRG6IkHR
7sss5lyfGICyAA0eZgbQzWB8M+spilHHHlFCpVrt9OWNapcZjXLTGGGIx9EW9j+T
Sqyv7aXEP6hMvzB3fmTJ1052/w5SQVSt7mn4RSizgoHYNAH9U1js0eze6y70kSBY
lxfkc6SjkLl6gjuIiPlPL+7wCF7fuwNgHu1D2GGcvtL2dxHDXuTf5qNPuv3aU0DA
sqzNuyIWufmsTNer5MRwzqep37OKWi2ogu1eVSWsKDcba4+GYBVAoWOmMX5OdJgJ
x1j9/Mbb2xrHsVxpQnhLORkXwYRf2Thpoy/1q923mJJM1MtbAl6wYZXmoRPIqgbv
RT2mraeW11aql/nh3JaX+RQEeRKO2+xReYZPA1idZR0FCsHvcr9s8hRlmg/djhgf
cA7UrbUG9rRmHaQX0wAc5aQlIb8SfFsC9uXzHDQwDtOHzj1wrvev/8yvQiWfakUg
pykIHcxuZAP4yjQx3rBeNDFSy1QYUtKo5pnrxpAP5dkYfpuknolSZ78V0lk8om0+
e7NDCzaVe85srr7uVrnrs+rXpJZjyJfscrwybT4oyWjN1soVtFiENmykVL35MENK
jGLmS3VhU2tfnzQkUjcL4UZeqsgrSYTwhO4ZnVN85l/EhItEIq2vS+zbXkK3hKfn
Wi8uN/xwq583O8egpF7smXDDpPyChwr+/Yq3HpBmzrmMs4fq7KkS+x1nQf1IxfT8
Px6h2wazffN+16Navnw88PEoKOVsdLCle/tQAQUH+vzC9GIhLJCBfX0JjJnLNENv
KggjMW60Oi9GBTrEIF6ux+3MfL5Tk8IyK3iaGC2us/M6vcYXOaSFA9D9xZgsl/n7
ZV5m6vzBF95Gx3C6LceyRKcaUsz2zvLuK9kid9SL3wbJTjSw0e+B5YTvN7z+97q9
vVETlyeGbO8If6zQt0Yf3nIm0l6kE08Fc8AMXU74BYJaQLEE8RBX9sRa2PufSBHM
VUU2rpFwp8WbkYluEXzTaqUaq8n+47P+4hEKwQIUc52dsYrNNrPkbICK68E8kda/
w7t0MzQUN5ONxhIUrO9am2YucTqyivr8OtT7BzKmGUqp+RvoRX6olj6u3LyQTVxp
NhNJxW6QcHE9BiToJZAZWFQLtVRxsaD4piLSGvJPRViHtaoQH7y8fW7h1rsesvfy
NCCkghYjFp2dZBXjVXvJYzwl5S0C2x6Ug2Ns1Ym6f65i5Uwb0Vm5Q6QeqPkPkTWg
e+wBo7IkN3NQO3H2dbXIt+HOD8BJgz5dvH7urGYFvUrDFNG/71kNRT0XoDiHM4iR
kwEZUEurMpuiDa+bcMtcLtifUdMrhb6novbIff4YTMeJnOCva34E13DIsJHZd5Ae
2Ch9TykSmF85Yu4+EXQSEyIQM6GeUQ/YOYNdnZdRQ7AQcnL24V5h3swwyqGvUwwK
gYiKYeYP5kkGcToleXrREwVYKNmvA7eWRe9bX0yI1zhEB0euX7YmSRl7WssqD+44
O7OrxQu44rYwy+gJvf2kjvJCrxIfuQCO1oNyYBjzUobVZ47U+eMRVuZOKON+KmcP
ObjdNFDTCoPHytoLSUarM323HsHJpvYd/Nms8dq1s38aFn2cK3jjIo6nHEdqWeWQ
pxDQ+a/Hn/1fc/a4GHZV0718PIxGrGPQiBc5zsk7g9mT0xOpEHqHsxu+H3zofFom
Egeyxy6A9VlVihjit+1yk0KRENpZ992orciZcnMafNSXcKwV2bNbQk/tmuiTRcOE
qmZOGPGehy2tjYdtdGNW9m3J0vwn44UrADF2T7Yl2XB/nmgUKjD81RQMO7iWYpoq
IJfyQApShP/zU4MZWJxEsozG6c7i1JxMJv6P9+9Y+GUTdmNGhxXuaQC3dnI1+jIu
+1TTM7mOfK1Yal8GLxxANkqY+cLP5xMJD8hZsj0pI2mgZhcx8aU6Viu6A01I6CiQ
usxxxl6csXfwLhN1Iwu0d1YXNml9sxpG+mSTsoAmbRISw32iW2oB199GnteMiOX4
JB2HtEmndGKBnuGfymgW+BibMygqAe8amt91iyX/8Jt/RcDmuS3vW8H49Er3PhWv
3jBwHFiUugM0nbDGqp4MZw8CqsgdfQvqqoMm9zr7V1LEH1Pndb4Zw5TAoxGmprmJ
/rNxXEN/HG3u3UVbzpoRhuvxIXHTFFgnhPPF0q9TujOLjdV5Xfh2KdiGYZ2gaA7P
7DiwiFynPMMNHxk9yUgt/wszZwOec10UAoo6RyuKyyxVQ3tCUNQpNhHPfrSluNR/
yRQb+tGT4vzEvGD772bAe+5mx8EL78VSX24SibspN8KE9rDtC77SB5UGHAMfiW7i
IL0j+r+YhvYJtT1/YVetciRSR7yFg5or3hrHNjMKuv/bqTrwwh6aOjPnO0HE3H1K
ZwMD0twsBB3Xt4uhMylQd63BuKr7ILYdaDUCFBCIbKb8d9Lns3R2uQwOjfVm+FAI
h+68/GYpKI8aSQKbBHCgoXjN9ZCd1EhjSozysxDes1Q5zPT0uXXLZKFTjWRCN7sx
CI8y9j2/0X2ZhtjaxfzvfqNpZ6767M3qcVvTEDMbWSRGf5Qk6M93B1y4SCmnlnRT
AerV5cUN7E9syLJ8KiQPZC7A/4pHMFhwoQlpZeBR4ZgQ3g9t/bRgFmGXiJfmcYHz
ktz6amNYlYtiVzX6MjQbu3kL3CkGAOEE+c6ViFRYthToYndtlAUxxp7k2itv4gaa
rF9XlTOHq1IZyzRGa/+psfQe/e3He3+83gKVOH6xbxu1kooOepz0w1kRoH8FwUDm
EnoM8Nzoj7ubAjqwdkyLjh6tRR6BK+WVLfmmrpd/IIV2oqjhxoNu1Z/S3c7Qo7lB
oyksl33Q/eAmlN8Nd7LxsMUX/+gtE/Ik5aSltqDaaoW+S+1RLxF9CJeAYgce1rL6
nC246VkcDpkMvt7l4DzD/f5pID7uh17jS8/qyhHRqz01+zylWEf0JB1X0xQa1cVK
1K6JGTby2mh2q+qjWuDB+e8NfMNpfhqDF04MtxMsWsJdovS6Go/iniFTHgioZOyq
njF6ImXYezeYNP6MrymgIAdu/GeTa5ZzXqtict9LWAAyKWUyOk/Cclr9oYRVeS2u
JuPwjZ1FQR7U3hUp+adQkO3MSuP7y4ER+YpZFzsR1L5w0HPQmEKOh779ZvsAB8wC
E+hUhYkV34/T+7lSxnxvNsC1osV28s8B+PmmjgaJnlICz98eSt3fa3s4XEdvqGdx
wBd694oY1xS2NENU0zvpxyJvn32UYRkbtfXZbsRpZcQHBzhtzn6VfjBmkPFcQq7p
imsGR+xm0P8ZZr/6k8gv95x2t+5l2Hj6ceguQjtD2BYAPwcBuvH5BPHYSP05qNlX
QZHi2pShmrLZNsNXXEJgm45TnfTYizLH31GMN+DJy5135vGX65LlQVRD+zP/IEPb
DY9ZtseS8kX4kyA6XFF75udfiIvqjKIoa3zI25ThduesFM+LHXwe04LJ6Z15slq2
OnSTEtvyYGcmWE9RfMoM2v1AD/8L5gHGtyRbij4oP6qSoRpF4a1IGkaBQds626lv
KI6ASvSOFnSq6kHkdyS6yIL23nRSeADdOsyk3jGxyGADKArW/Vdbd5Wdse3DEJz1
S7kWqpM/GZHNmLsRM87hokPY1bZZXVe8pmirycUk/zuqIVQa0HvZjrdv9YWYfb1B
Dx6sj7HAFl5EiPQ3SSbvtRn5wiN+4fNLj4oEsScyUmX7gDDs/SBPt3SsfBj3LqsU
jtaDhXFntXBvN1Z6oiJrb4l7FtA8zZBSW4hSK+davQWw2lwz7C2kuft3qoUtj+/+
lLptXJFQqKqDc5wJ5LjrETzfOOUDaIXDprtgsVHd7fFhFr34UgBFyDc3++bcvVwt
D0BhNBMNYvAM0guW7LTaLpf+P2SZZVPmGhRg5huHAg7Gb0oDLIbBCwWzxAsqcnCv
0cAcrP4u2z50qV91zPZvJzv3KpSW0k9XZQIgEyBrbxC0QAPi11xXPOEeMDxK8eJ7
V1o/KHsnICyfUs92HydQ4AKHM7cjzku75xriCuOsAEOZJ05mA/eZM8kiqVoAvbz6
bVvifXAHO/K3dzbcC+MSHU4qDwz4xMddF+eAyYl2O4+q81VbCk/nyxhPL/A0suSU
o8L0XE11giiv7flT+oLdVeDmNZUOBP1jY7yRUCFnTAheCvOFRadtjvYCy69LG2F9
XchTOJClZ7YMvqqYrGGHkTQrxHoANMXgtfIGKetSz4Y1+BhzQYY0ip5YvinCqWdk
bawqUdhvUHeHYO95Q5C53eScqrP1Se+kjiXiQSKakBagaRPrKUQDAEQOWYU/VCNA
BAKUxC1j1BxX2YVXTN7iK6X16a2pdX9tOs5X9+j1zknzlt9vMVrOtRm+Ys98b+dj
qdhOnpMrx8bp+YNXWJyk+BYC6gUh9ZZFFu7T9PMtWJxO+f3YZgn8iqDInfcXQR++
M/aAnzuOaecBUh1xdQXmmohvnMqfgpecBHJ6ZjQU+p8EqNuJJrBgCrJk7T2Ca9Ka
lZYfiQwIEsoPbe9eIBIXb0ZL9Uy7IMOntAXzHlb7+7aX6H1N4Jgu5vv7wLiOLJtC
YJ2axr21MWuNMi4UNnnhTcNuFqJwpBWbT4WuLi26EI3z5c7SWbHkP2sCBumqiF91
li19gYu9Fol4/GV0tYVrN+eF6EBBjM2GMjTpuQGcHhR0jq85rxJgZXaBsAscpgol
9+wY0xKM/5v9g/mXBXcpTQm7WBA5Btw59veN5CDTbkEGyKjjaguh/JzAWWI1yIGj
7tx+dCjeXQ0e0Nt1+cpZpW5OGYMcWIAdS/6h53zm/FCxNZtB/DVebRz+fKUHyjcW
h1MgpXX0R5JTRwzNCYh6RpRhdKPYSL+cUBF2DEXhCPtPysn2H7YkhrExKRQkMPeo
Oz/Xg794n0kVf+GzPVW6JrRzgsDFFqXlx9zUNNRvas5Yj2k+PmRi4rcshW8FbR8f
RCBIoq9n2B4AAlN28TyHr4Gmv1MYVtS6IWXAlZfSn6fUZnK7dST+lG0rBkMUtgLR
qQzOCZaM5b7p6IWLi8ydg6l6C8VCp1ec6ksTF6jjPCoSYepe4Nos1tZJCtJOyodo
YF655Ip1Y+GYiTwJCyfneAIyHbIiLFqxRGkNjARBpXingBFfjPd2psFI+6PUa6tA
5d9TN9yBTM4ka74ZfcevzbWfYSUBGgF/zneQbazSaP8CR7AQ27uQrLyZVk7GG0El
tCvpryR0e4WDDX7yeKHsGe54t7FfXZOBhcYBUdE/eSe9Tlv0PLMIgvUFT8VI6jaO
mVTdlhvdlz9JmSUH7LxGjT/KAO9Bcl+glsqyIsaNRzDDOJWGmQ/3zbz2tZNK5DBg
uz5ndG1T3zG24J9OoqCCD/Wt66oc4eI6zLNgUh2AjHdZaiLuZsgRNT0HE83NkIQ4
EZZKJ5RqLbiGuF4XG49y7R1hcymCIDlQozXBOYGIe9Cu0ghpv/9OJztHamNNqo+S
Cu9LkLn9SCUieYbGvO33WfvB96ZzXSi0sO7yTKSxXMrO5cHtXimLWk8aXCb5z8sv
5SpC1lQ+3hO2NThata7EdmoUJpI655ya49vp91qj3WXDnnC0MjD8i4RFW6R1rHn0
87ZdUrCiyvZRZWn0PeQi9h4k0vvv0yRVoC3j4TtgjRhJ3oViWIf4nFTlxNx8EAIc
1dH+mtdGynpRAD/6ZXOYxjrPsD6d1wT8K17xokqbm2bKJIuv3OfQ7hGeqqkk/QYD
y5z47utGJVVDUTnT8u+/zxHTQoDNloRhx6bBm2ZsiVOUOfoXWAEc0/y7swQJzx2a
D7PxWZ5g/t1WDTOTMJWFP09+YhD2l4h0rcOdryiaX0FRzhM9E19y1fBF9IcmyEbp
ZnRbVB2V6RzLdFryqTh/F5QXdTHAS1oYqRbGHLYqbYmj4pwDf1GWgkDMWaNhaWvY
w7/G14DllUgc8ggzCFLD89SvhpeYxdrm9vf1gEHzeo8MWP4laoSVClP5iTHOwXNG
Ge8meH2ZtK42GLMIH6fcq1BvQPoOdmSbbmIM5oPUFEDJv66ZtqDRI1AWBVWoKnV7
O0zhJwDYpQUj3xL5He8An6CdBvR5Pg0/LuGuyYBsVfgDJeTMZYWVOhPMb09Hxc9k
WQ47Yt2yCSCmuV9sZrdbGH1zfTu5GpGlC6ImXSmlyY3/QdQ+4mgLjQR5UQIVc3Lp
83CXcZ06Q6FgZ4RwkyliuRO5hXMUJPW5Y5riX+X26R6fUgdaphJbIFPIfq3JPzFb
TV/nJa2da8w/ndGYEGbnPm6th7R1I0kCC10OTdLk63r+xueBdAAPcXQTDuH8gwCt
uDc55nh6+pFteN5+5XU6GxnHugoeW3MwS0bkjAbj/kmSUNKsWRusy0+sBpzNRRTe
AeMLipsMTaIqUGnQEc6oHes/oo7xXleJ1UEeWzEVIFzMiYV+O5oVXwnpeKLPc6HK
oejMn9rkkADgg0QEYYZXZkwr5vcIYPnwA7qTVxqXNRetRqykOBw9e7pzQwSwEIaK
asrQkP0HAxkZiHMaDkgzTnNyjKUFaWwOR8591J9I/g4Seah1KpgCj2IQa2+5/ei9
v52o9KDjERvE7OJUpbj5WD/PC5Ny5QAZ4QUzB/qMfuOXmoE2HTBGGQJlJ7YZBKx7
9bDi5k0bZNS4dnCt8yD6IvPLOkx9dWNGdFWWZqlpz7fn+oHu1v7Px2SrdHSBBbuJ
0g7ab+6PEjN0Dbwtjpi+KWMyoxvDMyIBspK/XykPGA9Pj134GJ+4+IfByxbqQAAf
cBn8+Ty0X75nrGoNMHK+twglYKkqS1HUCUAAn/SxDQlmPSfbamhVr0OSV3fVicqO
TdRG4w2g5YtqGaTF8eLI0nnquGkGSaTu2OrgAUuYXYeS27CtO4svxxDAYq3dwMHc
q+MPonWm8wY+gOFcL+zwcsxLClwWRI4RYijnzy8ecmFJTOsi01UF7kNc5R7MTZw1
Z2WEdZxP9QXLWa/E4jjywSqCAdiLgNXwy5yel/OgjmxSZ7Rj+DtYPxB3LKa0r+Ew
58oXpKEl5lBmnGHlJewjyzZBFIXygBbua2RH+09rZNIIyPfH0RpOle/jKWw7Dh5H
p2StsyRzK+R6KsfzIS6MmTFinNG4zXBiZPAhFUfOnn+8yPCLxy5PNIkfCbcWOsxZ
UL6gtZ4FQ1quvD0PxMU+ljpx/buNRjfE/aqLFP3ux7zHmOM+pEmvLSr5Wl9/eXCh
papGK8D3gYFoQzPy8GxPiHIDpV+XB9b+qxxOONGDI0e6L/9pQ5la94uDpAsc2sou
XEc60vQBBSfJ2KMMsB5UZM5gMI0r0VUDQdsAB+SDe7PEtDNMXzGoWTiFaSYyfMn1
hG9kpEs1OVcVtLBTtr3sZY4sECM0B+jq4cGUdgonpmDm56oyEC6UD4E1EHmg2JbL
dEmyy20UtTl6CkydUUiDDTm0X5X3ohNpk/DZAzUDoUNAlhIOD9KdpVCnuOK38WeN
bp2lgIX6wEWxMqZX1Ty9XcnM2iMP+1/l8rKqL64udsWSoW2nUasfZwQWImShVoov
DCGTbT6wuCunIDtocDDAuePtng8kNQh2CJxTSbQlIDboP5GyahxFM9Srx1RPp0Jd
Q/a4SxUhXA3QCuReiceoDp/XspfKdmDst0jWuiQr2c7xwGnijfUX/LikiV6OLMzD
qjwn4YkxH/w3s8A9M/WVDpcI6UCd5yV3XQVKa9oZiF0gQjg6uQoWUL4SVqU3B4l+
/hhNUtLCFZ4PmhVQ5mTv/LSRxTx5R1d1qzcxhmdAPEQipgxrrQ+sUgiAajZR1pBs
0ytkvGt8nHDW3/56lC+VgRRnKwmKfpbDBQpnCYigq7VGUx61VfMMti6KKd9/UInp
llp/AAasjiB6fZBejZwBuUV8w5MOvpUkWfKFEgZd6N0hHLhPGJCImuPFvQO9m4a7
Jgm5RaoeG2mig2mUBW+GsD40ud/7Hjmeu8m0Fbr+Zqf3wRj2OOrAfIkmGhrJe6O4
DLESXZ1+JeL5OuazNzGcKsyOFSH3EcmxIZT9rqR4MHAwHrFzvCHrEhK17+O6g09J
oDaKl4muvjIn3jBYP0dhTInSizQYa5A9+exPuQs7Ft7kbHtW7avUvnUEhCxJFrqL
HNFKbchOnzmktaXG7A5ZTj9IKBhqx7CPZs7xjw52bcva/yGI0R4d/B3LLS11Er6K
XUz60swG1Pj9v7Ej2YFZ8YwrJpIUpuu/QGSlPSWjV63bvW5N7RSEhWgJT7NJGihj
cVBOo64ELFK7Akh4WDEsHlI/7WPhUlvVTfSaY9WQ33PAM9ze+6ndkFFjf4VQeDKr
sD6z9wZPFFk7kw7tR8T6b8UA/Dnyp3p01R14o/IlP3tEa+1YZCWls6+Lj+vQkArb
aYDd0ciQUsCYHzL8b17tkq3hrZVZRLpwWD2KwL6xmgI9nwtJF3jCADUu6DoGhlXW
fV4hkbBYQmvLmbotKU0MBaho07XNnyUHxyAyfTctokPXMmoZrzmrtzkE3GFqgtPi
87XEQIVTwaWIzRQa7Cf3osYU0lXvzwUQ7mPDzF2hIihpx1dqL6cHiA7SRmd6Yu6s
ELv7uQWrW/jW4Vw91PRzUDRYyr2WiA5C82s/SLJMBkLosj8v8zfbmXI4995vqGD5
XYRc+aLME0JSoAndMHOC81DxkyVdAJzvKZ9hq7e6s0NwoUQyR8Im8muuuq2reuCg
62Ne11+Tm5E5wBfncXn6JHaDam/zEobQCYqViGzegNo1Yzpq1vSX+NzZRzzN/Owj
Cd3zcy1LaoI3qDNI66vxEoIYl3iTVaa0g49ORpB97Z8Z9E8WrSKF3/ZQVfICiDd9
Jx/+qLN8m4xj79cSkpA0dNiqASF4lGEoMLBhPqp/LPMIFylpECZpdLsVWQH2hh9g
0wf0jW9sUujkRFzWI2hZ+zHOJER5SkfZDsdddmdqRXgGRzBWEYORxLj9UaBStCyq
sRxPRDOAF7GGIT0FhQeeet8YPguMGQqqjVrkqydQdugSTcVqo9KFn2WG9L7LXUNz
wtbsx50DKnk76eN9DA/4kdVCrQOtjijqXzvR7xrEmVIPDqNMMEcGns7gvYiawfnN
gsqyABDxhDezzkorYmRTcU9UQk+tyeJ2kk+PEHTtyTYxxOlgv86Yo6RcSExdmIiu
QUWTuSrD7gCGlH5tTmRzipcQSsm099vtLkNavHFTx8diLZ8mDtZJlcjUOseWrgai
FcokXvMxjEOgp7k0Tj5lzrJXhDX7ohEu6rLWz71zNMlniexfJ0WmxQ8jzkNyXETS
nGE4bQ8s82ZhyoxlSqZ7i0QYcTBYyfYW0Q9m0fJredjxeS5uAFVgChuThFpyNVfZ
P/d18EcrwBXhhdl9+7SgLj3I8K8ZwIp2+7OJ3E21frhywpG+pQG7Vul2o1QGd7eC
u2Sk1AkBzXjXkW0VdPX9GBqfMqi7NULnpDTJK0X+j4k6xl9kZBwjY6J9jbH7bETO
TXJH2O29qoqXPQ5ZqQHtWiWmq49xUI/28zXhyNxdfr+aH+JsGuSlfiMAVtUmfTRW
ITMOrlDNOVE1B25Vx46gcDIzeI/OAsp3QZAhqBDAW+8tdZz9vByY0uY+bSKAjDFb
+K44H8gBlt/flTuMNtIB7CPBf4mPYPodZVvHz58YGfEtPZZ2RAI51slFSspsp4G0
MG51AM/twZA7+TvGRY+8QsLmutES3XtZtCeP81Lryn5H8FL70zw+hlgyB1R2WY7y
nHa+PxtQ3TFykdoxLQDzTGO1GlFx1rw91KmZK6PltEilGCoamKnDHq4nXGToLROb
7Bd51plL37spblWSv4j5xQELVHM6jYLEQfFwTJzj5EIvyNstoA3hpMt+uNirZzj5
OX9GBxH16892nYl0Q4vlRTs7sy7Qjs2H3+1KARnd8CHX6MnYJZl/pYmQcuThN7Ya
lS/9/CUvxaRwixkNjABXHR6NljSUP3d1OV42FNX7UjtHLDv7aTcHUrij76ev/rMW
BeXrnGfHaYDHraNG5uw9chmF/5obD7h0ddEh/wgD817jq2AYgZ8k7vqjeIEAiiNL
GLo8UhH7U0FjOGdBaG5A0Dl5YR/RUQ6Y9PQA934UYk7LfDiHT7ltgH3OsyFSjj+w
kQN0l0OsHwgPSwfuX7u4OWlD5M/adRJj0o/riu2ND4YsIodNdQ+KXaSXxnPTanQk
KHyppB6TEnJHD1F1nXyCdBPSslI1MZA/Hz8ULBnWNgjmZs62V5+erpNBABw4y1mt
1xtEe77yrMoeJeEaF+Sl0fy+CIn4PROgWbv9XZxqo4suWQtEcAwrix8cKgEIkYgq
nb44/2BRJdXhwcPQNUZY2k0BqAdNRg0wPCIYpNrRENG4LW+KvJLIIZo3hwvCBOnv
V8WnluVDVSsV/F1qcgoFuvan7OvFcuIbUPcURhWRMKGVRVvjPkgT5afntdYYLlo3
65kddfGvgfi57llYXJa73ycpmMG2VQ2RE3FMB1pTM67XyF8twzgNBtJhwOjIaig9
RGAxpahy47IsstRq/S8YnK3EX624l0Nz47c1xwBLzie+wra4Jtw6b1kjpt0lUd2F
Exhaoeu8u9sLwoVtEO4DNnjZOr0uYWCDqyOTWgx1gZ5CXIbc7q/6VfFzbsps1jDS
x433/RdxL9fLv0cFKSRa6EFvQIUC7HhI4JZAAgasP2+dZsdn0GGwOreveTUqe6pE
6cfxGR74Fc9Yuwn9tu74hKkqzDbJ7GVr2Dgu3IPLCJiKVStRarqAWNrc3ecaJqjB
ygm0Z9LairUNAFP3j1HedWbiM0nFdi/sMNBYgL48bDzOhQ9sWRGbCxF3K3yxvw2U
ZipuE/TEDLFb4ytrVS4csq6ihiOYMLSFw28IruoqI0nSiCLUluzO2kxun64ExdFW
JxdIyb3FxsGGU22F3LKq7npaaGoxy/vfJikuutfo2ERgUl6DAQYhDcHwexUnf6gm
us75GcekHSNB5ePkRJe5qsPurnzD2435A01XrpaWPWjKgifAPmZrEwFa3LPQ9Vn+
jUC372mAxU0mHkAFDDL/KV0VEq1ulIZrBFxOst7jIPVmrazEb4EUnVVrRE0Q9u2J
TO7agTlu1iSlxHdPSz0qv/lJxI33tSGmSE4frhr760D447CD/NgZdDsjK1aStvNU
4hVWO3HnStmaVwIriOLuyxg6Mmm9u2RmMLs7RGTgJgqbMiDpkzaDX3RuVUEs9EdW
Q8de0Xb/RajP22H//g4/t+/H2bxi2NMSdMUnEf7Pqyc2kqk8kCxgO5IiQi1MIWWX
hZB408mzzPlrRcZPwm3ZZ8L2vkahcBMoz1j28ly3Hn2UyuKoY1GfLq7r/Y7MCed+
28+TPp1ozaDiwfW5hgImEhUwn/OTOWG0Lil3WBIj/EkDVvEU7a8ZbCETN9H/UntG
Zxd6ZB/lbp2Y3+xnkmSOrZmFvx1zjQDP6yLdPvzd6yycCI4oQoBBD1KYcF/O2vv/
yuWKl6cAeK02f65zLGd0hUP5QhQ9W4dI2x1Fdndkvqz52Tnv9awXXkQdXmh3eEUv
67CF9haXtv5NKjwoM84LU2dEwZPVXEnkiWSIePVaMWvqQkYP1iMvp6hhaMPDMl7d
u8j7B2heTqw51L0sYMtEDGazFW0qdpSJirhwg+pM3iYDFISQJ+KfciIK5m8BopQf
9rjDqQdiAAJbzj1+tvfdOVMPGFG58b03Xs8vZfq9IdGb5FH5KCV43TdyQAA3QVJa
6vXAiL05O7bqbR8ooc8VkdWseEhLvKHzytkpFYFyr0Y5mGn6cmXlQqDCJB8fWVwE
nd8eTZRzEPyLXI/PK5fAPEwWDw3VP7gTpdx0fzPlMmhM/gHT5eb628olpcNmteQn
V6Be7cKgFVUcG0Se6pz5ke7Fjrf8S2Kkp5z4Sl88yAQX0hStuZ8B96TbmXDD0Drg
8SHaMSl0+AVEXpGZ19mTRepn5Jv8iHRLowiDWtUzRjzFtyKRscB2sKcIkDl52me6
e9miBHLACBAxN52u+svViik04B9T/l6wvqfqhEJjTcZJr/mqYdHPIye/gdubYJ8s
fKnNEcnwpM5yjaHHqkJvaGqVOgwMCqbSSHgnGz56yvabRnmiOeiCfWd1Cf2csi1P
m8NpXb/c3zMddze5bpUrGfplUa3rAhwj/QgP8ONMXR3r9rIanv3QuY4m+d7oq+SG
oLz0rqd4og/iW2r6hvg/gbcQKUfpYEban21wccrW1y1Y+V9D8qCLD6bnfLZo/NJD
goTTRA76BymJH+8GqfsZ8Cs0RfmeWdexxNPtUcH1fdrI8EUoz0+oxA84oPSd1EtO
camgTwMV2L9dEaPTw0lVBkFlP/nrDXXNzwSb/cF0C0meqcybZ9PnbcXTGUKNDXwc
dGgIArwhn6e3oPOzaPOcK/YRP8dBtok1LbZnH00Xo42LzqiX+1o7P+2B3w/0xtSe
RHiMTHzxbTl2UZiNHdh2JOxWd0DFBniWQ7irGhgFtRLcXR61zU6mHYctw1ZNK+iE
IFcDDyOrHksQEhJhZxutFSVh7ddBjyVxgIbqK2liih64V5Gz/mY5ARAcq+DfD+SW
uNSWWFX6YBtgLHx9MrJGRz8d5Y9pm7Ckg6qNWtlyumjerCFEXImekjIIjf2k/RDJ
8QLUs1KkIm51yp7STALZy9xgMhwzvktVZLVkry5SKqOyCOtUD9ROCR9VQE2eXjNJ
GlQWKX0I8QKoj3+ZuvpX005l+BEY+wYKtHVTrfkNbxPCd4UbyhmSdANDFXTjBtW5
D96QIluWn8tP6IVL48JVeHOe++INrIGWl6WwFD14sOSkL1+Sg/Z2AMrsJGqAWXg5
gcNC7DopVH8DNUMvWTRLxL89euH7SHrYkn5fTCO7ESeiKe1MUGl4AmypEoj8W8ni
7XQJQGBLZk3QftqRwQrK4hGC1NxQLEd987HeSNiP210IT0tG1Rp0A+8rFwj19JID
ZXShNe4lL/GxBpBxNwG78BO7nFva/bDMYqzZCf/WWJlXPvxjvgYYCtsukZBt7EDx
Mx0HMJ+aNbVRTjFgC3zpsYXb9L7aWlffoELCp/gZRMcQ0eB/5Q3tmiLBU3G2EgwW
WRapChWePAtl+Yi1Zrn12iuQc50gM+V+T2iW0Jqv+lldey/gLmCom9BotXQf7YN+
4kmx2M4aLJD9uxjZlx0jV+SPCEQOwBXDmtFzgiz1yVc2NxdqxiOosNIcMiipnehz
TkB1gjm75DHsQOolK4xX5rsEIdsUnJpTmXRkjd5gT5oyH0LjlAevZjESecmpyPOq
wohHLgdeeFbxqSQUC7BFR8Yf9p2kwQ1WQGg486vECCsOYgynAtNWnsKRjKr3ni/3
pcrDCju/2vveW0ZQVltGmkTbln3ggs1X1EfqW5Kc0BZi708M0lnLTDkZqqDPv/KL
1bi3bkqsnjmiErKBnrmQlpjy3g76ENwavujSUsZ41tejo/oU1lvHy6bXW/lRbV8K
72KqJvfGzeltx9Kgudl+V+F9WtEw5uOcYT4WiqQgeZuXA0m2IOJ5DRFZKRaJZpIC
ikCLA9qdQZzfqmSc7kVTGxSBvXanG0MOFa0WixP7fX9O1BtvOz3jFqPETp5faARV
0y0pT9CCXAiNtBswOHRgooNB8UWTCNeHMyK/JxAZT4gHtS1sKRV+V1PeYCz4QL1k
HVukCZJFmQGb6SrAYdbSk6P1Qg2optDH/EYPfNumPSzyKJc+8GfpGUEOBRRnoU8P
GBGralI62WBdDlJK51b8HGd48mEsFuuh2S7TYzgS5yYpd5Hkaal6hvnvMKvUhNKC
jDGfZ7TJKxjBQRNNkAXhOSEltk2ysz/iQrECFHby4leWBy8aEGxqLvaz2M4zRsCp
hklstHwULN0v9a2r03S+G03s8a+LuT9pqQ2HE4KRkuoqHm7RbyVQnVL08vuO+Tig
yooR5RBuyWgfx4fXo45G+lg8PaOJmv6RXg5MfHR728D9QzK8DwCbyxthiaIU/+gO
/ukqAD3KwQa6Vem7xHEj/ydLRPRszZHfXxmdh1gre2uzF9biml6GP5L2utFJ1nA0
2VfD3xgXQuvJhsqhovpZW+hpJlSOfiOIS8P65SuXXRrfoC8uAy6zuNE17VoauZxa
/1sixdpJdXQR5kQklcJcWVg3XFZJ0mkuAADbj4IaHV0N9YYSLHO2/gXHtqrAYT0u
naYgVZw3nF6g0VQPSH2tqhnEWl11ZHkZYri/IJ/QzjBMb8C/4r1lE43M95IROZm2
2NY0EFSRlnL7tP9X9botqfES7iqC6NK1EuQuWKozh4QdiFvQfbWUMMsbLFrnJ8fY
jW2dKPELLBTkeC1Am531hl61HJbsWbdzo53PpP7hW3f10i4X1Kv5k/fY9uvE56nK
5jVDbKJfoahy6O8Fn2+RwDWLAtzxjk3ApBbDlhyauIFH81KhX4QsXUvPS0co8+op
bpYxSc4I8N9BiZkpAPm9EO6O6BEZMZ2A5lyXSzJJeiRRNTTJDJtbrSla+3aNd5Xl
gK4zZMprSZOXY3lzQCjb/2dhEtn4VS/8vqUGaJGey9RII9J4W3zrGCuMv+ScNTSl
CNTA5ykFkkxXjOUWsnkxigxDciWGGdL5Kqn/mkwFvLgwfbtPAz0v3ZoUbfM911Qa
wQYgc9xQ3dg/xnF+xYVkBItdqdbbTbPSUukazaGammQlq+6dOzT+6yiMT85FO1nF
IB2489Ax/7Jk22xaSVhdAIasBNYqlhNS+yYtwwqxr3tTestQCyTSG3BP+T722IgL
Mlppem0bQjeQkGxdzMX6zRk4rWtgz8FSTHTykAeV77wk7GUzJcum/VAp4KThYowQ
83KltH1V1r2A+YR9WoZmgJLVJhOLAoL5r3aACdCsPheKadZ1qTqtiLdHg6UtGZEj
ASGdVPh+ef3mMUfwkCRDyN+m8N9OpOwaKIyfEWEJ/KsglALhqfDygCNm96YKHwzo
DmRCjnuTGFHTS1C4EUnuKvtQrANK0A2lA9BVL7NHWy9vA0HBggfqf235u2VKSV3u
yPM0FZVn/QUip1dUvOobjuPS3aKMoX+gD69+AVoGGp0sI1KWeeOAgwjqbIPqxo9C
lhONzirDK5AK5lOPkW8cc10Tf5rUeVCcvAR/KwgJ/5nh6qSwxotTRJ38rJVUst1w
oZwl1PJeazKhhi7oN8opqIRYf8VvswarkeTQHz5iP6Pp2sAlUZvxhcHz3L0pnhzJ
+2vuMM65VRlzLp8DzcGkSsifCgnkxAuswEizHhfL8TffuhQvQOlb00gQh686v66f
yhFp20kW0ul+Z1QM1vy/QlhbxUs0Jv2mxhHY5mvHPSQPlOxMrYhOEvGJXG8+aN/2
TV7dOid/ZLiwZ4I/BqlZM8W+iKwViH5mehZpce/h8sfyf+YXxKw/OFChqbhX0VEr
CTsHzg1BF2lI3Xep6Jgf5OxedzWVGfdo4cDdQ93uKtz/KVkbhSdkRxp4xSEExu3g
vI+St5o3h92/RNRN8GEustERUUCabtbhHd13j9T+/dTKj0Ml8JMxNYMrBgr/V3DZ
zkzCPjDCsMCDyqzyudMDDwI0HRNLfki5rOxI/hlPtr5UIl8NeRKMKcgq2kfiIJ0K
pgFXyrlnGCI9LWfqgFjyGOoZ4fDpdGNlApqR9Qg79Zj90vbeCfB7ZuAMLcDLcG/A
uO0dsESU6HVFU5ukpfCAJ05kRnlHIehLCiIzKB7kfW0jqhn2RFT7+IDp2ZSKvmWE
KA2bmLPfSTXkdFwHLlFCjaGPb1PjZudjRfh0j3INBtwfbvN5BbhcrcVacF7qpMlQ
0qJM+B2uGYjsqQQT7STBMU4B24frMLKGh+j8yc3zi9p7RVPAPX3VuCZWjA7ixJSD
rqkwrdVpHIaNbXrCjt1Uh8TCI8PTn/s12PMYQKEnMGKBlQF5cavmiu7eOImpsqs1
tqGGDY2HIQ9J/yNZBE5ZaI2WRSHu1YjxEPGLO+JmrRGl++ziQF2ouh9f7XtPj2uV
1qlv+M1wr6UN/jWkFepxE5MXkbs49euxTZ4vC22wQ/+PRuFc7TRODPXT7cV/pyd7
uTgPR4z7M2OmJZ4ZOUGiA5uff9UjsemTVQwEerAPCAGYIMB8U4YK1XegztMHi/i8
9LWGYTHTHkiTUQ1lE8nTyO8eLTbVrnepWdtQJOsVZtDazReBXgmb1cgljhL32d9I
vWk1sxeFhzTXNn7BlxA72JlG0+X6LV/xxSuMiAB2NUj5rhFiVtvtsFebRv7kE0pe
P1JrX1ByMZjG/FxxTigu8Mz8WWTpIeb0+/SH4X9qJY10jFatAUhfHO45alcJerlT
8GV06xoWONHM0F3NB9vaFie9YoMZfFFSWciB7yoQWsdmqk5UROcITbo4OXnOePzX
EeTBCN0Kj3DXqAy0Cljup8x43BXQoWxbocRGaybIj7CFve5859blpdKehT6mKrAm
oSz6che3UV40tdYUOkQH9ikz5eDSCpvpg3oZQNMfPZ6LgCowyR7o5lo0dICe48w2
+nyivokeBUW16H30myj/7OOYyorCBkZy2dZdOZ05KGb2XnuBRkzRRBJXBlN3mbgO
OtmE0vVUl8aV+VesdVPnjvb6AVvOXxm05rcs5UncesOnUEG3Ws2RxPIQDLEPZIa2
Bk0TavjrVuPngdord5cTE/MFRX+gaWgxs6ao28yUS7ZECrUTmfQ0o5pdkgdh1oOg
WISys+soepJF5QNZtXHg0ddaGRj3cMJH62f543LigH0iIypZyoZwLVdACUJx8L6F
iMgeIrx+MssG49VFoQDRo8W7hyRYbcPerppD8f6sGsmXiOd9sRqEavUyRiVt6z9q
FDvnRxixkAtxp3TGRtekJG/NLpK1WgB4OR/kRwl0P0Wr6JQMdtl0GsRamdcx8L3R
bbw08gG27MuVn/KVJUSVJwizD6bMxPAZ2yy8+UI9VOF9bXBqJanxetqDZKshqgMk
73jxxo5W2q7qaYSZdln2B5I914HUyLRm0uvwm473LqfhkFiOJ1Ptvt3xrH36ALeu
c68tUKcm0yT08UuwfDV4NkL/3g+oFj1lFLqORlEcdVcNInjQtevizxDQh7KPkex1
1ITLtR+O4z4yxvlfW7E/j6vWJv2kR4XeJT9H5K0Tpxd4sf5/a1Nr088E/hDXxUvr
XNwtXRE6H7KaOL2wQ1ol7HihNvCX0XhdMsNxVCvonkwgBW3rikMee+g/GQ9He8B/
ecvylp1exX67U91odw5/ercdkkHXS8YLjdWDSd4Nx7B4THN/0KZ2oRkVmSy5ihFa
RXBb1BdlJg7fu2pukJNqgPwFfWF6Hm6bWuLEcGN55/4blPowefpL3JxJ3RZ9TYvk
cp0rc9UcYDCf16wE4N4W5HoPOXq9GyfMJPzR0NA5E8gcY0vSWXmwRp0H7DDzGDet
yUn9vCt5lZ6gfR8ReDDJNoWGQS5RI4UuEZAoyMQLfDAhA5bHJOE4I1qfAC9vaIt6
6W+j8dk58N0XmspmFBTbTOcbhsYdTExrZJb/L/mmiuk8OBpjd3iwckmk0csFcKGt
mo2Y2rbWN2OV8y8lN+6JIQ==
`protect end_protected
