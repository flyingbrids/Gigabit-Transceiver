`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
HsDLwKKpUDVD8pvrDi98QB/0vmPkgNu/GrrXxCP9pb286Ln8k2JV7Cw6+2p+PXSk
ZmYPknHxHzdAtYxGqE2oxiQFGVmCLIjWrcFV6IIDoJmgR9bAiZDAH2jnwQ1d2bYa
y1/+NfJcS34qNejBOVI3pm7vFnTuvYMh6M5yK377dEir1P8hBN3Kcg4f6AjSjJWo
pXerAjOxKzORpjf37UZT0bKXqNlHtvtwHiHYlAPwvAwRfA+uNOfmDyVj1h7KYd/s
d7kFdvlR4OgU3BzNLJbSax9Dql95kWhN2fqWlNw9yOR58aaVbtp5jznGfQo9YMRj
10L81Ft5zFsmJ3xaqxlOEA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
fwehLcp0h1mxbnbboefI5dTm6INvRaI+kccf14fcFg0JlOoIz8orN0RZ8ovWIUIi
Cd9jB9d4m4FLk4eWf/xVMgzxktJ5rnBi3O6fJqFk/9repqQ/s+WKRUy8Bx7ZE0QQ
oA6O6k31hckhMI2lc3n0ny20abs4gGcfY4Q7AfvJTao=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10912 )
`protect data_block
FUg7xShsUu947bPIPZlYpzRNdWpmIO1YWpTOClyPIndPk4fFMHxdSKdwJ8qG3fPu
YLz5VWdFZj7FR7y7ck+BOzccdBU3NdJvuYSH2IL3YLYxibYjZtXUL+ytKBSoEIxl
RpYb4yndMKT9Wb758Ca/qlEwdYxRp2h8JI+7Cj0aA5S0Av6T8n/hbksgDWYXVYNe
j5YEhV7Ehk3YVQ0Egumguw9qzI7ft23DyQ6YjIMjxyqBFJ2JZGQh0l8vo/3O2Z+S
gtlN61pvWOgHEDFmRp5M+xJD2bp9oU8t3kNCmGpjKRkameTOvQ9uYqY4bXy3fDu5
WGbbGVdvMzhTT34ocrei+S0hjD4Nx9TMofs2madUbPDic5ALbo07NNPSIVOYdsXJ
2WflwxINOlUIwtjNCxG42X7imaMBtlUss3sbv0WEcyCawRyYX1d+dAXZ5Cj/a/JR
fHTf7Ge8cHDrYI56VbFNX1doV4Uu1J84QIJyZpZCufGt4hqKSloMuYYH/ixj2JLy
kp9ZPU1c0+AIyZIwew5/yM2YkqpXCA/oPMbAhm1UAVonYG8VCPjAd5/bARxXu4A1
3kpO9q45BC9yxwUR97EfqGxxMmwd4PYkLjP7RK21vTvlbzW6r/WoYXh+4I1IlAg3
l7gSD/FoVwFIkb3mCch2C8+uW1ii+ELTp7zDL9qB5uSPJtgCUrtv3MpTpq7fLccq
EypEwZxfGLp8KHDFVHxHOyMsdRmFjsYwjr32sDbH2Aq5JGmmtgg+rtO1m0jT62j+
oYE3eKUzk9Cs0QYU+8LaIZpuqq6WW+M+6ALT5KnN5uN6r+lUIa+yfI3LnwxCSrJE
Kb94mkH4aQ1fWHOCvUt4WSfm8ikzx29eLyCNYJkvzzRMM9QWGSMFAb1pFktxpbRo
EScaBe8pvNt0wWjqinYNW36jH+s9TncT8nhfdJWfDivn63xEogov1PmfnHP/QBSk
e+cl+/nQ8h5rhgYPhlrOxODhNX964RtOc23nvrWAZviKwSqe1+3VzQJDwdQRPLND
ayn0w+aWNskg054IfC7/GiN2CYNUiAYxLT75Yee28HbhF5nlfQQTJwz4XalO8A4v
UvHjMQkfZyHOOKcLnS/SYsVC+xeCXYKA2Pv4W/16UBF6AqK1pVM5L9bsAvGcXUah
8yDNdAkK9u3VnXd8yBj+MpJ830T/jKsnSsOVb51cLYyZg/uXu7gb0RYWfl20W7qK
bdjDSMQFFmjZSM9mtfsdHobKRS1/l/gKQdqkXKPU1kO/Ray5ahKG/VUxqUl0buda
/R06P2x766wuCtPK/xoanmnUWtljLFN29ot3jExH91eXQ4rjrXpUVcYPGXY9O2gr
HehoCnXKBZavkLoO6aslmzjZKo/+PCRxbj1KhOQniXOHegQE/yr6aMcz8VmPIEln
aarGk+9WDpeLS4y4w8cWEkz3CN2trJuigSB4MOH+/etasKyYfsWfmajGcaCwiwsJ
iznyOItblSRtb87Rhe4LsUHBtW5aZ6nyS+OR3nenKJIScA34mx6SflIPCm5dJPog
/HWDYOsvjPHMmGg4QTBAVo+plERo7Owu/Pqome4VQ8mgK31zgMetcGRjjA//st15
TVrNQ+8WWjyl2gkXZUfJDlB1dB8jL/H/UZO4OvqNJxkdLC8vyACeeIsdZkh6tJzK
Buv7bfCgeRMIFWuZG0U3ArKDEg5K7Ppna/3egtC8cs6J3Z7VVQrNpTjLUmAh+0kn
C+Xw4FH6wCZWNmyZ5n594n4fAxItkC8DvwpLJbw+fFXfhOxhBb/+h9Lb9LKsRtiU
D3KCZ5tf60gkNywnVkqOBBIhP22PU4UYGnRhDP5U++lZ1JKPB620MMfsUGA4HsCS
PSWYakMleWn7LIDIbivCKNxCniYDzohtTEL+krMj/25Z1fM94Rf7jcx6qwTxHMGl
32YKQGp+hqnNaxsIn9sfyBmh6J6GDSjv4OYpwzepczbPH/T+ecKIRWP7YjVC+F0F
SVaZOjW5JSmYbF+f7RjQOSnDjouu7f914QUKZytm1LwS7d4gNNoeaciKYt0FSu39
tG85aXcRhEB11aIJEau44iiaAmlvF8Rvgy2bVvyuuJT/ZCXyldocmf6r+ZxQSVEt
LUpXaP4HVYg4nQrGWltuscUNDs/vhl13QSRQ9bhKb9S+nq826Nv/u0PP0+hHv4x2
UGfCt5r4AtLoaU6BNybn1j4wu7zKRTVXNi5VTMu6aoZu+H0sY8+cfDI9srA/YhjS
8YMWyqc2m/I1ZUyotDvwQAjXx5q/ygvtgpxMOUunlxR62zEM3WCF3zL2Xg+ZUcRh
N0ITg4TBRwrbm4cWDYyx5IO/jUUeNavlXdEFlZCtCr8hmRHrqAyI7VNK+bIL4n09
tNGVGLPG7phJb84d4T40Q5xK424W3z8nZDDSPZdzq/qKgtdTQY35repXjzMdRS+6
aaP25ZoEdKI3jRulYRwF410jPIwJUlJFC2xk9zIGX002jRi5a/HpfRFPm7Ie1du8
FkIB2dl5P/WAewQs0PEqY2P4yGTTfxOMYClUmEJOPN151b7hNZ9OVcGX2NSUk0wG
rXaJMFewPx+LXJIg7hw2WE9S166SjcvtO5m8odSFh0+zzt1ypC/OpXB3q9Ykfn5n
ggrQYGOWHQbV8ufGb1ShMScyddVWxXJqULoVRAii+8a0M59RME9dvBNpFJCzoK2l
H/P+rIllGeYuR9opAdHx3hlCAttxldttOJPj15/rYYqpdXZ6RCEuhOxZgRPgUBz3
/BQi8Ekv3GB85VHXOqH0xCO0FoP2+GIx1GX4mZxpRCtMbweJBZHOv2oDoda9qF1s
GlxeasxwuQe4OPXaRUmVYyEPHiq5A+CjJANe2SiJAY0V8GIUnzdNDEblQ6EnFa+c
qiH6/daiw8wAMlAqnwOLCini/WGwMQi1Ha+2IRM4pp6FEJS86tTxCmaMo6Czilpo
Hbvta29B9i+V5bDfD1kUknG4/dmOpLmSH0MQlo0jT8fNxMAMfhSaQUMFnMCXynn+
t6X/Ycpgt77VNdj56gDDy8OWTR1StatJ5KJI9zQJtx0ObJYv66Sl9CLFjVoJwVYb
1cOKDsdhJ/XtBpn9judmFd7ltubpAJpyz3Ro0z6zFDmYyUSaXeULLMXHEUIaahVL
4Rzh05hlBoYTuBGC8Pu0kLD4Xa5xVkxVQAWAtdwTkD4wesUNLUJSSlBrnWQn8pJZ
9k6qKcZA9i0vNIAtxZFpVR/+fctc+QniSxzpiaP9UTCWntH+a6gHH2sftJuA394i
/cJVtzsotelZ34FnqBlMgjv5doeWVmY5cbJUE+qVGAaWPrhfAIJB4t42ce1hRogr
M4UiTqZa6Q24MEHpebsXYL+Rlz5fPuSG6DVUuA+0I7Uqk+cxRKLGLTzR3EDOCvhg
shdB6wGFZF/G+wi9yu1H7GPyyrfHq+O2YJMvW3tiEWwixtZcBkWoXXwnwfCNT2fR
FEDpyd/eLf//FIvDJOHn+AiVfONRTJTT6rB/XTDSuxZonZxCLwX7v/lhyaDVHrZ2
UDj8H//8R5A3TZB6xkhjN2FEvgo/rC9lW0Esbgk0nOyODuDxbulhHKPn2rT5tmwU
01rWMc6RG9+J6/P3L5YIb+d3r+ti18QN4ZeAACwsZnSx4Z+zZ8LtOm1frBSuSkMD
bgeHPcwJqWJ8JGtJ0cE51tkKAnUjKwGBGGs4PYv9adX9+qdvnxMsbu0AYv6N7uVO
upGo3dcv82vZVump51+0VsbQ8BJTTxhJYjARC1V37PTPOz99jHMl/FfAex7f7uTm
BstwFPDOM5JyZhcEPDhOkT3Bo3P9MON/AmEN6z/4rg3gB7xZFM19mSMEvyhb9Lc+
GY/u/Y4eUCUuBBjyz2VWaJB39vhsWVjUwXWQPh6VDlQAvH7EgpjoE6DoqV2DZ1pk
48+MrECMF/O4plWt0nMlO1kl+JVSWkRiTfiIx+EXSZlnrNRRNX9zQwcptvs3Ta1C
d43bAGsqSobgRPmwsbtyexQPxQsnZkRuz1sdMvuaIKSKKvR0vMjx3QZrCPjn6ep5
Dy8fCJv0t2YtsF8fnEsrGYxuUTv2Wxy6cqY9KbIyRBWVfUSwklHl7FFHlWoiH+3N
6aKkZ9W0ha820WEkJ5L8a7jAOf55x78wJJQEviurfj75mJLD3/MZy1VUMY9RpXsE
690TenNsJmkc4pKacV8J88CUDgNduZfV/9KfAX3FnPzJBL1cDUE+DneNTL18IM2x
+jFgfZXqOPEk322+WmdEMBDmdYzN/MD9tHHVTDj6Yyx4u9+hxkXhVJJpNmQWNPMW
n3upubqfzI/gqkE8aVh8HuOmMh2MwljHTyMTl9FwTBdxQRP9tJJsDJ3SNNH7hsWx
Xn1xjsxkr0eSzrfe3oJH3jdBz3jS7Cj1BLZXFirdQdG7HCxMPHZlCfkmBly7H2ye
/KZlMI7X7QV6w3gLuNb3JCLps3ODOBUK96ZoF3KUswc2/8PKK/orasFFNjcNWrWD
xMxeiWoValIQCmGmq1sLla/5DP/7LQOQJJllNASibD7mZlua5VFuxKbkeu6NsNVv
Al5JZy4Z0xVH78Y9tdPZLPGLgw5cP8lPT37bXJ2fb0IBl0cpiSsGbw5PvRmXhdna
8sE7Rwh9zyuBNCfOexuoLds815WjYFW765N33MAzWW6C39Ip4YUiODh6kmi1HPAO
bZthWssjbfVda5eBZxGtUTFKh3/+WXh8lWJ26rySGC3cTmFYsn0aByHZv046D1sY
Wf1JLUipeOW8M5VsyI/Z/md1Az7rEgbBfJ1dKVNCwcTCjxMGbOCJWoAP3a95yM5m
99AD3bnECmcXGgwvjZbySIAZaJyxtBX+1IqZd1udF2roKwRW+K6QhwRNpRMkgJw5
phMQR4AUuiat60LUY2CpW6witK464BSfaoyX3w77QNLUEf0jrunG0Stbz+JnSd/V
kM7SjmhBSP3UlvQinCRoIx4BuK3qIYJURTn5PDyXf3SQJg4Gply3e3MbRPm1SQNw
LGxkFbFRGgS5aezMqXgn3HG7UCf2HkQsUdOX0kMc7zHfmcHrTwqJF4doeE+wIJSX
DQZbPJMaflaHBVtlvHWdNH3OTIOUM0xKFazGHjSFZp3p8vYgGsl8Mogl+f2ANx0C
23wcs+xpvB/0t0i5yDswGzA/VQAgSixFiMxTGjSm98yuN2FHxw91yUWSsG9o9g64
LV2BwxV8O+7SALfPavACGT2MDJ7hXDq9JC3Gf5qB661bcyC7fb8e66jDcC04yyB1
SDLYjEed7oUifAgkl+uklq/0vCQuuyssZeXmRtszc2MAKvCZTkrIRnJfGqh5jyQ0
bGUJ/91DlE5H5ADxuWAUwTckKOHoiv7RycSsVEuE9XSvmdClRXV7F/t5Jys4sg1g
Cto2rD6G+ztTGXs9pE9plPgc9ndRbL5200o8GoVjwEbqa/EtXDL0L7g9Nu99KTkQ
0ITiVIE76djQSEtGduZEqfOkEmM1vym/SWT9Ex9PgWiMs9aMDqRVaFoWDlomRQJm
O/2lpPYd+Zl3mYld62FsZFvHVFC5tze0eZYVZwf2ShLua8s/KIZsBpgQzdEq+yGp
SHSH+4ug/XrrB6uw7TMmMYNlosEWwakSltV7JG++8prAumecK3L+of9MSYDfIlFm
MA5woC7Ux0eMuxEX++axQZ9NCNmePeuj6DGheek2iJu7bgkwxbsJSYQgvXL7RwCl
e0YUbPymDgIZGtnJjds6jg7W5LSWcDvgy6wM24D40aJEywJlfZw82wRGNP3QF6Jl
Al5RnedUWVnlJqOlJPOcZsOZ7GyzqX3YqyTDwEfRs91TCmjqUf+zrtigY3/oLZ33
rew0PvL4yHo2lf4ZpiucrBsr7YncXibRXnz9qJUxlzXM5z9BHdk1LimzPVV0gHDz
7Bfp0Gh3yNyPLcVhdUqGl3pAn3aeXuXPvPxFrmCa/pEVctCb7uUeXSD4Dz6YSfkl
IQXrlVl7ufigtaSW33KsUvZRVphqnfYFzm/rqG5a5c4L6RC0pv1TPB7+ehHcXU9h
6vauqkn2OwQcw/OmqKwC0ELJPD03daEYbBLQuYHw09fDvmKovWs9Xzbpcy1WoM4N
4RjDnwSLgtyfKhlUX6SnHlWu7F/GiizaHnaaDNZf02yAIrYF82l6DaOVLBqrW22O
JJu4oDJc212J5mgV/wqucGeq8v7Mme6/aR9vqY2eDV74ROgrw0RI/WR+ow20Jimk
LyJRjgUoxdkKewXL9luQ+0lKepryFaTwQ6hIgcZCWo711Bns3VLjh49rjisx2pkn
po2wUr2qIIeG/WeYWJY60kF4rVanI/yNdHe9mD47D3s/ZKQiFv7CeRwvJMTRyGQ4
VxrOJIR9w19dZ0mFBu/avBRJEjBbYMR6009uwQlr3V8dOuvXS8Ys/geis4xtfl/4
Af3eY0Ar7gmnvIFom/KQQL2kjxusRl5EPkZLg7FWHErBLuM9eDpZgrWzr18zKCml
4SaIyY7esTRuCh1DX/Cp/pdhjZsRQiBF99OyWNZFYMXcks6lwW2KfBcKDOZoVegq
MjdbP6A8p3C8uyKA6E4Zz/R6+HH8HFzIlct44k1ENr7GLEw/tnZFGMxO+5Jc1xEf
HhlcFYlzm3r6xtfjxT8coqfX3U8MnNJ0Hb97Gg4tSsAuduOMT/Q5TPUnmJE0i6zi
Pwo0kI/euQxhZNsOdF6GWju2ia0rWQGrYZjEofMvK+nydbZs8opjGMnAS/FsuX4J
WJwmHpkGUzGP0BJHmL951rfHTuL7JsBmcpPus9MORPyZHt0LC2tqi1yeFNoeDF4B
z+Uy4Bk157EzdVHtrR7ZjomESY2CrGP8EqnAbDqEqPp6ahxIzy+CUnHyybGH78Wm
zpKgVjJhCrTur4Y2GxMSorvbLadYS4Br2V0RmFo8EJuPKIPg8fCsDeY+Q7pXnyet
K0JYE4StnqSfY6pOduvs0WhYW+YzFYoS8qE9L6wz/nePykAzEWcHAV3gs6nGQH6j
HNPQUsBKym4JFfNcWHCCvwU3ZNdomExukbm9QXI/ogdMWDvIh9GQ2v/KzYhAzzaX
f+IwPfhfWt6ha5FfvcfHddYE+omXkbd6LdQRIWdB6a0Nzxdotr0D/ElONcSriZVI
iSjv0CQTF8ynA70iRWUVHrPA8B4Oc7naDiszUDk/OUFE/CPuGiMa3R5To5Z2NTaZ
CXwWFWgAtWOFiFprsBiUD9dlARD7DVyYXoGISNLrs0An6jGPWy3lpLUkz5WMyMz4
JwpWGYJWQwirOhEI9+Eh19td5YOZPILuHAGort8Q54mvFo0cU6F3cSJMmd3awtpX
labydOPBOlBP6cotrUVcRQCPxOHTd57gyj1i73P/D7BGqKHeU3zXAxa9M8ykk04U
EIEWza8fY66jFJqbhkg67lAIW4N9c3eh4YVSHKz+sATK+x9ThwK79MYEHr8VNM3j
cWqLlbhUk7C4/IFEi+QhSrVbQCSjshZ6Nc8Mq8QRQ1AiK2bSCjXWsT0mG6H8XWPk
59rh1FCF8C2UzN57v1sVya9qq06Odfr6BHEHCAe/mjzdwCb0V7+BVhgrm+tTpcmM
DRC4mpPqWV2DBcRplWQxB9YZja2X/xQfofqTTCR0yq36T0d8cC7YH1xsgNf5nUr+
jGSxp0dHt2G2980yQNTAXHx5sSXf+4g5LqjEvu/aNnPGvHF1wCorgpvqrRykz90C
5ZVrzCnf/i6sQ4biudQDvnImK6KZl0su8nWFZmLV9dZQzzCj7t7GpqnR2Z5qqyB6
JESugR7Shc3NhNcziRykOiRom5HhGUt3RXEdtD5ci4aGXK0pTSXTkcAnoFHh2EVz
2LrU4m2yy7WVIvPnqVCjZaUND9ZXvGuqie/DaM+ySURRf+9hJtCnPHKOKl+XawNH
a9dVoyFW/Ta/G1d/y0MuHHSx4ssg0ncOjT3bRDUNmlvXP+mR3BKaJr8oDobEPljm
7wS6+wRy/X3efv/t1Bn8kG6CcmEuPMFzt/7puwJi5mAeQgHOKy4RyvFnCkCCvRJP
+btMQ0HNsmbuIbSN4HL0iltLs+NkMD2t7Qqi31CpvZ/xJtVJyeh+/yeRL1CNDBmy
09oUowiF221Kr8FsYvoS9xB5Gb2HcvZShZW58dCn860Vzya1BjyaT40gsY2mu6Dt
iS+H6pJl05kH5ExHsMtC5AImWdbXhCJzJxbN7Sx5XwIKMRTP6lXT2rRqZvsyfkoQ
nxQ8Mmz7x4dQQCjLi/DmGmQA3GfQ0Ly4UBGU82HYvgBwMMMhkoVg1+gKpmIus6NZ
42ldKuBpH0B89EZ+22QS7MZxzQG5mgt2TFIG8FwLnzmORRQoVkj1H9o1hSGEDfIU
skiPC6BHNSHKfl7clmNBvzVVnx+mo1axmvFrbMWnZIaR7jMYUztLCgzaG+zlgwim
es4pqc8Xyv3akW/PkS6u2W/B08c2HJCIZ10viGZSeciME+pxff7cHPoMRviCS44j
fWTBFUbNsmHstXEVyvPYougBZpJ1L8SPg3AhCAU5ND2TXrE2hNiv1HqafIRs3MBS
1cJ61Cmhlm0bkO8GMnChNhQjEoIRhH8rMQxQjq1PUaNxUf79eNRodzSBig8rgITh
Bk793H+Ik8yqWawH5XpcQ41kC0c2RpPUTaLf7MJrXi07y2qzJpAjQHoH2ZmOGex7
T4Kj+CTTcCrPu5UhC4ODqiugH/Zrxchq/j7EhQB/yLqnsVp2VG5ynH94AFaKF4d1
2TwB+Yf9nbS+TlTCN9B4BOGI2Zc1M/lMNnt2cOIA+K/av+Ap3ui7omwKG47h6VWm
hJ5dhQs16puqH7+bFzoiFLWDkvCXZZAt2ywdpav7QvJ8Wsu3mOUg1XhNGWY8J9dl
kVLt+r2hD22zuXN355lq/r5qvcfH/sNLsIouSOuS3nisiO1clmL0+h6NNhodpnNi
yELrTcWjyUjkkZP2XiBeNWkz/yI6Tv28Wrg65yBI/GORwMr4B3nKFwUW4VUVYY5B
Fq6u21QXnVwGix6GsBmm101R/OyBfm4Jfy57FK87GwNnDRxWLJ629JgKswI50XMm
Ip3H78Nu+CJFwePclwm9YBvJTChjODddUfeBOTPt8Jb42J3RoGP6KWJL1d8pWEJd
wKJkb2x61V/ehmDid5OUg28RbVmiq7b88drIGiF5iioY1OVU58uD7WJB293Xqh4V
Gf3xPdNQouyYgwGfEp+6C4LfANbfx/0jIyGMa12mqNyFMfWC8hd7TGGNR9GUKhPX
s3toaykExtkPyHAEx5IGfWuE2oXYTjYsqkLO7kE6IKgmSWSKEvuE9Bv/j67QFKtT
QS56MTrPTqZKqlcB5Vof6BkT/vQFsbOZltchJiiFVWVQZv+e6g4VFL9svv2yDsHF
0f4MwJjfBXAREpCCmgvfeVjBBHPEHhnIvtc7ag7jpU4LgViCXC3GTKFDj7uC6ZPP
QmHAqMaM8wAALB9ch3gQfarmimaGkpF6ExSWmjV21cxBHNsor0wzavYlUF9rmN8Z
O/kbDIZp8FARUngGUQu6OY0LdA7qqn+YhX+bVkBZfJwEUg3S/vNXctMhoIxN1jcC
/qaoaPRgQ8q6W7qHkYZE+bY/pYBgNi4mcOp6DWVzE5Gmn0uvLrzyE/NZFTPvH8cj
vh2Eaj7QXm/eLA+a/Ber/ncZEJcYr3BIYSuZdWPidhw+1Qg9mAGxzg7fxFbTdg+y
7dPpM8n6oLtc8e2sbcerbYUsmHmViByd++mNwT8CR1Z6tV5WKeSZZcFPdbL1lbFz
h448jElCTQDSj15dMlkPPyVc4uHn+QToLUb6R5adItM3xn+TyBvjrcCBUeUsXk54
atYonE9isx9aPgi3t1Y5rINvSJqI8OPrOyV8p3e2Pcpqer3o14NB1oOJ5L5KsRH9
KRd1hAQNpn+0KWZ+mFq7IE3GC6xR6MmPQwyMQ9V1d8OKCT1MXJTkRqKD3Oaxnzn1
qEQbuhImWBIHC8I/GI7MpGggYCHRBw/sph0uaK6IN/azaHOFUTo4py5Ne2YRrS/S
eGMRa80S76C3IOh/mMhy05z3SM6ov+z4l8s5y0g2YKkAOCVVX3yjZlRycYowZ24r
yZjp6ATrbbpeqgfp+JuC+skthY9opXXlWzMnOSByj8Ggh/TIvXPan82Jo9HuDywz
UnwTOIQ6S/3LzzUOzI28N739kOtQh8Z7OlJy0s3vfSd+y9avnG5zaRzL9GPRmRe/
diZ/eNOt1GEyFsl8H1xcawvnJ59gz/HcxKchkEkkhZbPmGlJF/Y3rJJ4nKGcvXld
FmBYzhn/VnEvFHOxqznNGUZEe7xgKwqE4YKbzU5JFxA1M2q3yUP9qzaproV5++/2
DMfciMo2keH+g3SpUvcucFbZGMYGYMurgeNcBYtSMNCd8BfqMs7htMRn4B9X8fxz
V9I5EH4MPbN2lSTQACG3FI1URsPmMNbd+oxKpWonO+uMEV7PTSF4cNe1fBf9bPLT
P/FTLCJpbZ/y2vCzrprold+rFpD0GFLKZJWndQihPBENevX8pXVGxWcE2vKP7Sjg
gO/cDJPtdFvaRTuRg7jbVv3dc3oyLU0p4wqIAbxgghzC64obT/UV3hlcLFVBa/wE
+nCGUIGhPlG6QlmWxIfeUXN4d3+G4Y+uT5y9RftenmIspU0e8YdOs3my3ToCRjxR
KmUvQhO+/kxPeXsCKVUHiJtnTBjh7eYnJwkEHVKPm8wpafK7tbVUkNS3rNv09lUh
ZlfGeAosiaptj1GSUR7ftZQa6U63pMNKuzOU7LR19GHRa+mJHio+Oyr4LoV9PAZm
SSFvQ1bmIqlPArmQKjVvMpSEd5dnMg7jnXejLTfE0IfmQsiWXcerRRDc+hwdE41t
h5PBGnUr+E3YJcimEXELu5rnHq1IirUDjKT+FwRxUpRjzv0qpeDrN9G7ie4iVC1q
5c0gadvmXUlqK8i6qP/9JXfe5U8hpOJE8v7qixuGINHw/17ZT3x+2AILt0xIXrCb
THvD9rOWxEFfW7h0dbseUlvH2e4SyWIcuRhV2RGRwGMOdWpmJ3vjmjek5xtgzn9v
f2vK8T2jZ+WONDQADJrASIQf7CgmK1lfLOjA2AEWHSesQBlApMrPcAWaXVxktmyS
YUEn4RpxTHjr0udYfjzS+tNErMP+v5MQ00EfNPAfeDyZ+BnIdVDEkEIw/jXj1JAj
sR0O+sJ8xWJmSg6SZysiiexKOsXE58GUHNr/ry4Ygd4MJe1eDAWTQvutQGhyGygB
eFudaTdexPZwsRvaAGN4E8R2EFV4DdBdVRK6yAPrkHM5zpT4GANEbnFKyeLi+a+L
2Hvbr1G9092qToUtd9BqSoADyqe2pIJQ2N9HtEczqp94KXsDiAA9HadAMYsmiND8
YKYiCCHu2NrUxsnnMe1U0tDAEjHr1ilN/oshOon0tBjh0NbTfmL6o24D8ov/xUzB
4Qiu9DdA04Eje2YxzChvUru778WJxMpzLSycPkvKWqydRfyN/YlZ1W59Mqujpl3n
M7hnLtJ3kT5CohdPAXmMiFonDFncO4e3Lci+vp324GnGY9YEtTizcYtWb2uGb+3n
V/Cc6Gx9QbWb1DBSeMeDRFK9v+baxl0Oo/NMcDmM5xVlhXcWv5CwjI+9XOaHaY9A
xQ6+MI8wpwI/PiyLGQ5ubeOa6FTmJwJFTliRtsSqTaQwFagj7T8yy2r2hAn7y5rM
IbFyYcOYw1/mqAwZsa9IyRVtS9PgviDuelGV//EYzfZa3XaehqAZVA3rzFydH5kC
krNkxN1N6MqOxQWzZy4bHyptwmZM9RDy/PpRqqQCW+pXGbIIRJLHFRtaFwWgCInW
XaJ31EiBcrQONkwDhSfpgTR0F8yG3grZCjdWT7mI9qB5nZNBy04IUVu0piFNgVXP
eCQDrQr8QzozpdnL9mj512pbRzty/qUmY/yZ+TQHxHgzooQ4ymH6O7NGUVZyElfm
bfFFjqiUKQcB1cFNMO3k7WK9bIXGm6Mg1LEq5rJ4ef8/XCJhAjcIqTgQ4VaOkLq+
3T3+EaKvDJSptijdIs1JsY7RvBUcomogATFjmS7IPbmzhX5vG3OQvj47v3KGHEKn
8gUlQ/oqsdhbBu5cMEJX/my9IkWp9JT9N9SiYuX69AK761vXJiu3VxrJpFIQ8UQU
QpBaiYfwFmqjf47VkcODs+jTLkfLXdJwDn9Py5/t6OE0V/g7adIWqNw89CR6kdSH
cQ/CdgrkfG57Qr1mG+38r8h6808cEdtKyoS+nTKuEi2YH8/8Hgg2OcTKrBgZ97kp
1cvrzmv+9cu2fE1+kI77hVUX5EQYmGerxukRAtuN1y9rdjLb+P9Eo7vcfGTY5TTZ
KiSJmSHI8XoiMQZYSUy/Ub1Ysn+xnhBrJZQvUD7Jk2Isii/BYYSsjKLIcstdFB0V
KRYEz+SfvPndQawHpvyWgnkClpk+Yxlynb5gJyjEH1nJ9ajNaR3dJHC04xz6l29C
yC2JEzM1qm/Bqu6R/qZwFRrLkmxaty5wBezYtvMB6kT3f7tOqVBxfSUAfQbS6jjd
fNabp8Ot4NtBRJXfVGMWS0WsGWUi73uF+suXJTqzvcFUAaY1guSRVQTUavAAKPv4
452ylshnFfqIns08xbsJMRjZmTGk+BBxeTLm0e2jnr2vpf9pB2hqMAjbuWIY5SFC
sd2bNz3pG+KHFapE7R0dtH3p9ZcXqDyJ/Utfzr3r/1BacD+0MUrAoQJ5TKRy35Qy
1b6jCp4ZDwqzk89QG9+CpzTR1WWDkv7Fvmq6ZxDorn6Q5u6ygy51uXyWqNiagAjh
bijdzV4NVLFxHXs+MV48DUsBCxfLRq0tmBAt39eCBweyN9bfzT4625JDMGhbf2Bv
qIU9ws3VgGynZvI2vejnrR8Rc+yf+mwBwrT/ff046hGLLc1L5tciCaMWShWPFMaM
BRv8v1PZajWLeMYNfW/uLbSo34f01NvEpDTvDmBbJ3ofTo9UMiwQdPHa/U77vSat
3gCDuRf8gq6csUEBmJ3EcymYuAWecKl+MhRm3wLCZyVdFGvFPLBu3tZjye23T/ZZ
uRc1FoKJdhk+X7URuD5uHBEiEQ4i5P9dlpCs1KU0mhkTn8TjTL22mZOZ+W7qVlGJ
wCgUoZzibsB79qWVcUF3lhtJGq92JvLlZlatwLX2sq0XY0w4B2Uji5sSzVGivZrE
5w158v0Vd67iN3Hevfzw9y31dKrBHWT5gZSpd43FeOsA4xlSmdpH/ZpqAefYiFz8
lEV8QMlBXYVfw+2voXayndEFF85QUtJlRJYI0gn/wQLPxELGcPfocHei1acIJHnb
Bux4AOg64gYG6jGjncWpssUxbw6IBEItH53fXdPvBqvg4PAfjBr0czB8do9PY08v
q4+HY+669RSuOUbZUe7B1L2PTHGaEoxgfzVA9lMaJYHmmOKKaQXIKlKflH5tEfEa
H+hlO8VWRCfgw03MZq5gQoBBAc5NDfhM0G/HZa4LuX45tvyFOR2SMc3k6Ym18MIV
9QVUXxjq64y//sJjRoLPDMvYk1d0+jFXEBau+OADd2b0p1Iu7YT2lQ+Yb7W/BKoW
C/L2Ta8oJPkArlKBrgAbPh9PGMQJ2cpK6VDHedHTGkxNAvtJdeJi+UzeIn9kJnJU
qdXB47ulneuTAGbo39suGdWBeALN8yIG5KIjvMRHZ3fmhBzH0/MRHf92D4bKj/E3
ibJ+/oiSiCmT0PaUTq5Ahz8GsbpSRzE6Liyzh7PdavX7N/uaNVymja7RsWd+EN+N
1hPuJe/bOrdFV+B0/NJXyyRuc7dB/Btf28hoXXOQVEt16KupTSUqIHmXVMAeNRjn
qK/rZ3aImBxKm7mLCgqSid0hJleIwd/CU7WaTASTAkY+UMinRpBh6CXViow6lbYo
Ir8Ilze8c8jdpypr4+Y2kvmnacLBZuSDiJz85hml5Vv/i+4pG2QVn4HI0Jj/clvD
7jkjC7RR7ibb2KPVfg0rs/F2cH1me8wCLN1jk1OdtpsV4kvb4DH+2M9wjFv5i20b
WXkRmc1wy03aHOEHRp/DK0q2JAoRwB5GIGBTiIzZL+mY46CX+B98Lgxoj0hErmdZ
aJFQ3EmxGfXQDFipIORaDC3b9dE759boc6r9LacUlI+XU7N2OJqwgzftnGhFX5t0
Q5Bm3sMljFs/T9V5mR9871lDgXfRUh9TIVcRhR44Uhr4aM4wGegl++0ZUbvLdGkG
S7+ica6+k3GP7si9BAVxboHYWG5wSJIZmGPFqeksunBjz8QjYLvjmY8SzqiHScUz
i2ksCeWUSr5OMQu4/7T3u4uQIjFUoQuyKjeFH1/axiu3cbBmrxcV8GhduCstTz8g
SPN+bz6/6euzN1BbyB3SBsMdFdmYQzSNzSRwNY8qnocoPwvvCWDeHkLMN4+6QqCy
myNUAda7Zh4l6MdVDfUCapsQ6pTK/nJDqPt9gyaWpNmiCZhRfdnKS0WVP9xLeUTG
krpzR9N0BX6iimguzFEzmllFxiGt4ERP6kv01pmCs1IarA1+izLTsb9GxrYG/hlW
3dZ0/BZTQRASLtD6SGkKf36lTrOx3ZDQRCd9L1mTas6GB3Ar7crPH/IUYc/+hSae
kODeKneXpLpNpg7xBdaGeg==
`protect end_protected
