`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
NbchhUQo9EDriBoLV5j4BcJvJdbAw8GVO7gTFQ4zdmzh3s5p8dSTSYNrU9AVIsWR
KiCZT00Uab4NzS72Sw4X3OteGOPSY0up4RBkrYT1/ndlNXwfbPZcGeTatGpN/BrI
8Gd+wXByXo7pLHbbvKJp+moEY63AifEe0acdpuwgzsP/JyB71WP21X1ln4RlMWPY
uvAWymCuSv3MC2n/A3otqQsfrva9Ieb5jJVWaqb/r5UxTNmpEs7WrVWRXusflfkI
mdAmND4ZCDXeC9Sw0yWFjtRBb8bIczJ5pZyNOsmqBblWKvzhl0NtpPLq6C+D0pUm
h4QR5XkSi7c0erbCt9mC0w==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
V1Vbd0WmVYU3WQqP6IORQcJlbAhZXARCSoLyPCs5ChuLYekWlzLIu3J5Ii8iWGM4
BICeuDzZDDyp1gOZ0fyfX8pzRCHO3Wi28/ECqzQcavFj23FznHnOiD8Ep2VtSF8x
mCIPFsYqGd/XZVpCNvuaqvjNpyvdBAMl+z4+3fVYVcc=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5952 )
`protect data_block
ttIXKKCZnnQuHeDogcK9qKmu5pTzU6CoOIVu+nS9x0PwQabnZpmtx6RtyHVv/Kdv
9sqnZ9ETpHjFdGbfGeqtuO3zmHuxJy39vydbLslfVoILoh5tuvLpkH6dII6NJN9i
ldDIGm6X7NqdGlsHsALiQ3m8N1r4ZZPtVXbyd0dPuZfXXZhnCHOIfbyO6dpvXZp/
GJiSvY46Tl8XudLWt29OUVV685aqnCqFUAbJSY3u3n37sVfcoBz6L9mRmybc9EMb
281vFM+/KyH/cspTAapFJdcCKUCWDwQdr/UxM/7Evmo2i/z+yfid+jHjNuHwFRRu
JzIIpvi6ORg+9k4pxQkDs2REu25XQ1mgCfjSYCTuoQBUN6PgvWEsu5tE6JNUO5L5
wPUvrlMf/KROWZWEOSgnGAjuLftC23oFFEbM0BpjsFXuQca7XSiZq5pmKFTm2FWP
VfHNyZyaBsUJWX1JOY65ivRVNwQLYVK/U7+Ir0eVWxF0HFmBW/KHgYJe1a4P8yvQ
inx8ZKj6DmnKoqh6xHE3FUrYuet+vaTu0EAGmJedX+piegAOCUAuDHET7cd4ycfz
iF0EjQwrl3SQDtS+nrEpaNf9xGySjX1RvLCevssC+wUQnxmFIzuMjyA5P1pVkEGY
ZGlRJ/PLRkx370YSl2b0fkg8fIKa2k7Mm9VQVGFtWxXoOz9SdYfVsmvbyoG5mXML
KO8CWwrqfreJezIo8U7dMMLcWO/0qswBE9/t4bynP20NORfV8R4gCVvbx96oSCft
doVsm3j9pyEE7alo1DT8HMElZFmSNVyjI1F6bkT+dk/mkssCAhhsXpN+BZiyd9V0
v2ED4nzLPyIjyC0e5SnkuRdt8Egoh+tKNfHQp7AqD9j3EZcujRrw6DRQOnqY+o1Q
fuml67UEARKDkVBiF0JYngw/zRGp4jfoUtDkUwhldQ4D0Z/CKnP/dY17e7Ko8NfI
6iYpSa7n9Cd2pdxVM6NDCh3ngtqexgZBneYWsvEjE6gKYCRalDFxUjOGQWjuqUoy
WEBsgFNHZQLMkv8R69wQveZ5o7VkFu3zMCNvIM1n8MDZD64VcOn+YUcgg/7FsEqn
4BiqelMcfwFNQ6tXm0UopHAkJ1Z/SzQQneBXJnU8Fm5qs+Pqjwb7DtSSLsAniVRM
fYgVazPGXhIwebyYdAd4Put7TjHK0z2LpqOQXv0QfHq/VxgxLLqLhYDuyGuAFW+l
Sc49QLLSGg7iEww2x+/Tff7aBuhDYYrSRpsvtFHywBH4Z24XOH2wvYhJ7ymWqn7Q
fEfGi2PSnWspeaOQtQzR5/4tQAqidqzkD96PLFa/jAqrbycwTWRxVcGYCInb7Irr
MqXJNo8Rhs8msJVgehp7GK72gf2Ddvol8/jdC+Ee/syEMLUcxb+12dlROY9q1i64
dit5EhmmFi/hxgWdE8Sw464duZDHo/u54yw4vBHoy8+1mdYWfBVonX4Ugg01v3Io
lK4M+spCzLErGER11IxTyRpWitJuQJmbn7I0LtyxqPjutIBabX8z7z7OKwUPrHZ8
QuggKJ4jTmdaykCGRSvAxnoKf3oFv9Y1yU4p6g55MqdoJFiEndPoYOG27jIcGC/9
YxOOvlR5JEu5/lArrhji1b43K2a2ZNIXupEujfTVOgjEFkBusLUrRzcqvePLdDiN
O9bbs3cGSqzjOFFW0RGtIYM0sufDfBOYrKH31QLcOk/hq/DC0PdOSEF0KNcawfNR
PhMI7Yur+79ctW+FPeeIDamnwjMp93Q9Yuc7GK2Qx1OpCRB2szB+1k9/Osmze1jn
iuee7YsrT5vFRjH3g7YBnSZa7FdZwsRqy5QXSUN2tszMMzkh6dUuhhZqjoSrG8fy
hqn7S6ciVu9NsLr17oVSufSe4lBg+7+nJygpOQAsK3r/y5S+9jPJeK4tIB/hpkHh
vyiOdWWZHuZC7U6mnfI7xvkGCzbd7duh6oFwzMsQkDOJSN/iFL/HUnBJykQfUfS5
a9U81glslz3eaVawXmKgpWS+MYyUEbHGJPZlLSSooAmy7hCAnyHxbhtpz2V/jT0V
tulbAmrcxXczgTglioJ9wsesOyhfadEHCGBJD+YKJ9Tx2QKlQhXTCMoypm42u3W8
rLOFz7geqJV2tnNbkyw88dtV9R6io10qNwAZBQn592ef3+kdhpTP1fxfuPPAt7rI
om9LQGjfil3cbabU9nSBLln37aZgAg6taWdzLfOE1b5jYdASSb8A+ROaqVwCf8Wc
fi6bTYEy1KdWbo6jM7I7Jxc/akpXHjcVZ+jzDskCFM2vkC4Ys1hPlluAOwzyG2AQ
frsUZGFRpZ70PjnMTv+qybGOkdOarVQPe/LFggI/SBal7h1pBjscSauGXcs/F9A2
2glA7Ri7tqOz53brDJZ5hAanbxCF1e5KKAhdzEP7P4DcaMzzS9i0C0XFDqBrFOBe
aVF9Er7Z4K8/lorjquJAJRqnC7QkadFbE2Zbq3qtKBLzup46F9GxEF4Mryu4Bkyz
qDrUM8FaXixz7/p1Jf1T4uPAtE1LpDL1exT3DnZa3GXAqW4gWd5mBajrcjxq3wxm
8ZTB3bTWOZQCDcSX6RZ2buxi1Q9YUt/jCDljt9dLDO2BVfINUvSQyFVkPCAhiQtE
oav4XuqT7eR/arMOjSNkpdSj2Xy8VTUda9kQBMKnC0SfjL0/ikePbdMPuB058lsN
PPu3d1JU+twYyeVEANl9JaXsUaOI1cfCK5cpdjQYwPcQoEelNaUChf8e8aKC/c7G
Kyid4bODrkUqJ8T5vG0izF5z3DehAH+fe8q7g832rWUqKM3QC/3u1Tw1TNCWmA6U
I7UEta49SKUfp7uSN5ZhOb2pToRN93kl1tl7jP0iBGSksmPPJjzd6Iu9ymMXmj30
5T9hzHVN26GOGIWyXsnuLT3gucpy6zg9rU50k2fO4EauGoAOMA+tv9wB7jBtbSjz
FcymDUS7v+mA1NPrM/GzSYaLGqK6IPw/h4L5C5de0Bog/EP+BRRU2YnpW5RHd8Dg
zyuCBQ8QfUmovyB1/O8jAgezLzCmhsgxs6CDCjXz89evd+iXC3jBn2V0fnreTOur
DXYpQpJ2+UrFS0q1pM3RfD8TVaV7LSR8Cyyj2HHAkBkVIXhrw9XxOVi/t3xksFH4
xNOq2lY4pKmeVhfJTkaTQ6d74U73nzLR+cimuRGOBK6rl1zbLWuJNGQkn8tOFNOr
zltLfRf5FziegtBRtUDi4Hc+Wo3iVA/ERIZkrygON67Rt6VRFqTxxspCXFraVlA/
N2xIZ9g1TsCHmzjHEAN5sQm+//pyRRxnE4DNhdjfDHI5MFvrA5ENjVOnIOBqJmLO
p5O6ObtJ9FLOnpp4m6/CRzOe5dJji4fDcPZa+dvFh6AW4b2uNHTSvaJAVuSKMRVK
4vONXjqNrLuOXJaWG4he7/88h8WEglH050XtDufBj0+b9jAhbDFYhFPWUy/874fg
cFSYJhW9Cn3zCcGBfdtsA4RoWF8vydyBVKQzlHVVeQqphSnk5Ce96gQD92RTY546
dJNbXeM+aJ212VPIfFoXyMfryuSy+gml8WcZzk7uyy1+nG317NJEMtYyuMGu1MbB
CQKpYrHUomaWRFLYj5zx3rX5GsTYgtXZ/E+VYUBlQue4d1uGLgEzwgcZEa0fUSnG
ZTutk883SR+utAm5JZ28Li9Mbo8gYCZGjmQV3vrH+emy60HwQVgrhm0q8tU28iay
fSEz5+ooJnhtM17RGOdCVC2SUXFJaHXX+8Hb7RRw7+GPvois3oWydgWUYygtHGzO
GMj6Aty8M/q+xidKlKOcQ5cRj45mRyA8LjUgTOLObj/VnVBkLchJVR5Nz0BfkswQ
5GUPuucDwX1S/MH6/sq8SWWf6sYIjssb0bUQzT8bTwdF82iZ9uYiaLKdGhGz1LFA
dYDceSeSlwDyh6Pks3w6Cfv2yTQNagH7eDrahmFpmDQDRlxPAAOT8QOrcj3M0alY
87Tkn5tFpqvhhkjVefn4n7YPzxN8qRi2gEFhSehJal/tNt/O7izlZMW6hJoKZqE7
GL3hkCZtYH3lYQh/ygWJNImvgG+bHadTKMWamuTJtgWgUlF94HJ4NBVSwvKyESB2
ZVW3hJoM8syEMXMAiLAAPcdq9CzPQ9qjs8KOaWBc32S31F5QlB0OD6Mx1I795sIH
ZEvYC/aPvIwo003uQW4zLz2UzU0slScR9JWlkakwVc+SfCLo90A44Ov4KpAGFEK1
q521+xdFKWG+dqmzzDeIKf+CUHDFAAmuoO1Me2FZyx8vbqZ/w2ENeVSoE4a6k3tM
Hoo3S1soPicVDB7CyxmyiNGP0YIno8NWy+KS4pMilcaH0et/FZEDlhsy5blhmdUC
vVZqiNOSJqJl15bof7jfx+6vd9PDpyJFFMlIFr05q1zE7DKML1SHaT1g05vRZX1g
68+QqUZ+R/1791/immlBcskObWVbo3cWI9kXVkaTYD2+K7PHdgdWdV/OkkqP8fOL
Z3SXrtG/DZPqx4JhYDguI+S21Hkcj5L6VqXdsjvixiUjsGjmNUXtkP7eClfgV0XA
esfXGmoNG+nw6twe0HfYuCTNe4Cq5Koc+NxnXZi7XEUPuwcUKaHYBTpBpNoIOoYJ
GLTTQS9OUXyN2y81c++TgKqyBxUF2zfpkPfLf7p9itt1KhT+uiwWkc0Y3wD5waDj
G69T+0wtP+qCik77fO/QBBOpNE+yddxKLN43xUmJaZSQKZR5zM9BudHu5Z4lPd99
+fya+Urvh3in+7HeXzo/cnllr+pz2LYnuVg4IFWlnTbRqbHMdRcoiKA1pYS1nKhL
+mQ6hq1ucQmwe9o25WnxsGkYr5ESAP09usoc5eo7CuPrxlIfN7getDBzwm3SgdFH
hAbOpXi276+teMAdRE9kL/izQ/FO7Cltp0gsZWUqnqXrvSICeQE10aAqeyd8Dyhy
Ya59FhhhQRifsruq4i0CkFkpxZOTBBhIkGCmw8cCEOBw3amRTZPDeU+CbMtNhf6F
AVvb2o30Two2OkSe/tv69BMZDZFODHTB7Ea1M0dsaOjrtTpF+CnHg+zDsyJJttw5
UQx4vS0YXY2dZDMDEZtwzbI+vpKhUGEhxdAq9eUb8pzWiCYoq072ZTP1p2PaURyI
m82Bc7yJN3oMQ/Bz2dxWJphs9ebeZudtS2KrcQp86n8IQkVgJar6vm7fMgs/ph3B
JQR+iPrFRRObEpZ4EdPuGJ+afNYgD9KjG2uD7F8fG1zJeCYMKTysACdmAzEbZ8Mk
FZGAifPThhKwayQmntp8asP88o6PvJ/84RvdKOK8SJXXjHkbuNL7mroDVhALnzL/
TP94zKqwAaPM6Su5Tp+JwPerbzMbdReOcUifPs+UCntt43Qv26+UwV4FXJHUtxmt
us0VNAYAoaKMsWe0/U4/x0sYmMNTjNn700LIentLoJlQOtnLtGk/vhY4bYVtE/wq
932UJfFgPHe4AWwPRRjW5IzwCACwJcZ3tzmDFVDGlBrvOxvhUccnJW1y5JzokzIe
mPYmiqcjJevJA2lhjvztqYDzOZBBwFwJIsyXMCfdvVxPo38uEIAfwA+XbPpmMrdz
TMXtCHIAzgLMTzQ1edqCWheZGJcqOEBz8Bq8+PjnMpfOXaGzd9J3ovQVzMV92nzH
+wbZoQD4JmwDq8bPg0sDeQLUH6xHCZdJP2b1fHkgddIfAlZ3cBFFv7jNHfts4DMk
XBWhsP24DUug9HiRIfC2ojRuFQpzGVwmW6DzLzxuv2NJpx8BCm/mpq4KyC0PzrXW
gZus3y7HjNF8JRYTsvkGDQ3L3FmYGOGiBC1VF2racnRwKREDZKimo82U885ZnyPN
d9U490yC1/f0j05Ugo04LkXYLtt3zuF/lzak9dPlpDgsnzRf4Yw8amfkHYLtt3mD
PyWKGRZlvwl3QSan1xBYWdZpULaxoas0htgPZjbFIIcLjH5J4vNUakFdTiln5Fao
qgaO2Kar3uL2vHvPUZl5C5xaB9KucsJTlRyZqDR0xByNK7P7mD44EasKZjH1onKP
tGXnDWZ0SF/Klyoquve1+IVlBOHDsZBaEc/cO1cGWKDJJObz/oOX/jZxt7+e9Uoo
4AWVcCz155S9+yUGhUGMA70cSftP4vQwTI8LME7lzCuwFThTjessXRpLOnsGiTm3
eeOufqbb8rvgX0uSuZZCD6MJNePM0e4tBbarpiwP+cWLM0jU1xcCPmFeU1Nu2mre
ax5tEw+w5KFVcJBDBcLj6RLu2Ip7gRe6DzBHsrEQCpeeCZCapBAflhoo3EuhF2my
wlRA4IiSfcqmnUaSxkOSccCEpWjlx0wF0DpepmdzcQMjo8dQtXQDp+F32zCrsDIR
bMVx7Oi3d39PU2s7WclNYQzZJPh1dYDypUSt4qIm3fSTTTPLq+podpp53Ddzvvb+
8n1hgyOLqZCb+l5L+IcnuNIag+YLCgmQ+0Bi196zXxzGCnjvQep/DxiwCNp3g+3w
EHbUJOMa0wLG2zJDp5EgVjjp5sIsX6qjT9mbBW/tSYfF4yEsrcmemkJYQoyRahl7
S+7EE0Yc6YJJbaLT3XUav6Rum4YHlZgvCOVevIlsgX/jep8jpl0v0q5bFQgIYdZL
Zz9nvSmHgeLRy8ifraI+rVS4J0vhXydIOi9uGt8wPy1tBPzeXcFQI11feQb80CUO
kUtkW1wl1O/Gd27lwQdnGTN7DwtaCEDLHIknW0hfr6mffOx1FkeSt712XhtGn0GX
fjqyt1XcayF+Poja4FlKLe7BQxBubKaiKcGxDav72So60U6iFyt6F2rKv8lMMnu4
htEYRYiyseiI4pkTPd7RKIkXBi6ujnU6ikJnmADrRh4SrjrVzYmiDz2MzVSOtHbQ
D7oJiNLZMWOvfV0wDor6hdoOekHbtbteEbU/F9/flaEd8WM0UnF/wOYYBWdY979+
KSCIyRLdlmsBl81ZA+2lZojDp8YWDveSr7LRdI/7WQG7r69ZHflRY9pcIBpCckb0
+72/QObsXvpDb/CQTEE6cQZvVdcmNpUYzlJt+wmiNtvcv2NWVng6ccPwJLkixhAf
/n3Gq0g5waUxCGWslVuKYy9O+xRxgNjLFmFRr2QW5XXtymGxylHaIWLZZskilIGG
smSLdXnRzivgE9CLfGWEIS9SmxHTgrHj59hgHxy+yeyM9xT3hyxyXiosqExs9s15
j7gr8vHGpBUxsUZLzFLZyRJGwrMDDmr4mBhyOSMckMpSNuSxaVK2zW8wHqLetB/5
kfWehWqXwLeRKFhMjGNTLAblJflILuSICjpL+wIEDSQQnPp5R6J5sAAPVO/mTkOq
KxALTJuN1QZKrboffHvB/s9S61zI3O81Agl1KI0SI8um5g8W7/30KSLlvIC+K12k
MXbdxo8qfC2aun4tXa3d/FwBgLEKiDFql7Bw5N72IyxS3nuXuVMOsNZjkzvEPV3d
wPAD+YCApwcI2ihKdKtcSrxMSrcgr8H/sBZUX7QPzwJqRPQvqy4Rc+ZRxoFc34F2
Xzt1jR/QhqSTVEmLwgJCZ2XgqVtZIOU2HcnH5YsxpNYLbNboKW9j3jthj2/omw6u
NZscvc7QCmJiyEI6TdDyX1k4/09kjJZuf1fT+KenQ8Pu5PgR3nYN8p2hBnZ7uwrd
qVF2uup89lLjh/cnN4VQ56mzoWQ9NrVkTGOpUSsvG8gKcb7u5YG8wKpblhyo+5TK
xj9vxcuJjWrTB7p09Cdf1kOeSmgbG4G+ZFlOkrU2Jw8RHaWEC3TpJlieJrD7oxBB
1QaxqWlpay6mZqtcIw75/r92aruDZJGbCsV/oF0n+a41J7uSxKMYXBqxqcZlXTsi
+FJQ/Sim/yfNOsp3aJuvRaDn8pYcyox0wg3sYeqXeYbEi3XqX8KzxQC6JcdMTBu0
SVHvvvNYQLeKcPbilNhnB+UOSobwMlx4I4PrAf9uo5qtb5jzwJq4h2GWZHXdRU9j
`protect end_protected
