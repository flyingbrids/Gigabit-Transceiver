`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ezMjaOuvl8SvHKSwhY7hBfXahy2XXNaEznwlTnNMW17nRirce1dvJw0l0kpw5ohx
fPzWxg8FNd2oXCa49nUNL+2XMVNZ3tRPe70QGFZ0xWp/0aK2QpUMxVXbCDo2dF8E
T/Dobnvf9yfgKKycjTbko3XjeQ8Qn3387G574v1Se0diHZYCxohlTCWi7EGafI+j
6Lx6/0iva63H0S/ULkT29ymRfHDxWCtLxLkbknSdFkJ16/IQrYiyahAKza1BACbu
8UcVqKmwIuwu8xyzA5mZFjvYTuDxXXO6m/ta2wv6A8dZsBvjnzl+ZeY8NwRU9k3s
B7ccCecV5b47W5K+1qzp5w==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
np/GGr4K2SWr2SayisuFumM/BW00s3ukVpRDXYVaEdXcaaEa1elCf/I8RsAUFDb4
blMM/XB2+eulcZ0XRGbUHkHDO1skZuzk4rKid8exMCSmfA97sHy5n3fGk5bnQmNb
jLeOsVTAfIPr8WFpuLGCHKxrweI1MbbHiLT/Zy7u3Zs=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 32672 )
`protect data_block
IJxSBBHy03mawkfweJenv3yUbG2uX80LhNES/+dlUq2tev2tzwZ+69C1BJ97fTG4
7xIBzHUODzHkijkd6BsS4Us3o7Mgj9BBsAdww+E2yDq4cFE/rQ7PkITnGjn7C1Lr
YSIwg6E8qxdkicj1I9jE8YLg4gsYRGSeOScMMe7sGkt0zbOcymhJEWM23DDt/qRC
aSBR+6r5OwZhzPC4D6yiJjYyn9UPZU8YmPoia7fPNn+KV/xUTdFNDvKIrGr3XmJ9
9q3XB/G//SCIIQfZ6SKT0BiEVJfivW/DFdNYepy2OqJHQbpzGMwX8Njxe6Wc8B8Z
bgq6+q6Z0j2h5E2CvPK1gCMVOZr/LEfvYrQdu8NEtzS/zxEo36v4bbEPpt+37jvr
hnNhsDC7tMPA+Byszg+7+RC09ko+i39vQHXENCKSrdeIzAE6VqHhpCw9tknPmvnr
Re0zSjm/vo9RFhOn4NWW1epo/gve6nNFB2XVGwDp9mX18U2Of9yKw3Ko0szIIEP9
lxZs3b4B4qiOFGG85rvwDrIKei4bZIgfESQEyM+QEpMa8GCcrPH8Kd4kY1wqMYRx
Ksud5CYkEsF5IHXcvbopuAvowLi2x5hIeSW2jKEonxvKvI+L3fbu3Yfobjdpk7NB
cjiLibTLqR+cI1MusK7V82OEuPn65oYAjIBAdprYZQFCOCk+ujc/BkEmD12wDGay
2kqMmvZGQuAoqQft8ybJgr1794Np7DwRdsq10hZ2NTXaMG94G5S2HYjwfXlHUeE5
mjhnf5aOd4H480USHcozKvkFJ74dpEUi2EKbd3fsyt6gKxbSOGuU6Nst57aJeK0X
x16BeF6d1EdFF2n99G9FEnFfshsFYI5e8CZ3cPkjH4wd9fBuJg7DAkeio8D/Ob2+
WySqmGK0sf3h5z8mXeT9XZCvaGe3Z62iXCgCSR1eXN4zVJgdtY0TQZ1mTLC85Kpm
LMrYCIxXGxUveDTPQ64503qIz+hEONf+KBQ+At/dnTXCsaQY9gzl4IMFpYeYSGOo
K2J+ddYdvD3geZdTJvrxWRCQJx70NxVr0t0HxU3wSKq/ljRgdJXetZZsCybJDdxk
00SopgEXk5mWImRFKBOk9Vqss6l1jgoTxxljOvnCh0HtTIM+J4OKcJffoME7vRcj
NWn0EzP0jbkenAjdVjEDus1nmAKlTq53DVRMc5GwJzGu8WcSeHZ4hNQwStR7ZTZD
TGduWQvfFsEV42L8mTfi19hSv2gvoIrR8TgIKwHdo+y9BnwFCEfJoCRoWgk9IDny
66p72C53/lEgWYGY7UZtw8Y76LnOgiHTbyOr8DEc2uiDn4V80duGfQJhPpVJP1xu
WEBkpSk+jcKlRvhvr4jqoaGP/QeNvnn/cwm1+pnccV6Bg2x6AN/O36t2GFNwGC8b
5Jv/fi/CDB4Z/CfRjGGk8X+Brg283k3TyBbZnz9rZPrlDHRbM6gj5eAe8vdV85MT
BQG0+0+9+B4+N/l8RH87w2xZhKY9vDmtY0mJbbYkWrMllZJOxL1bZO1c1V1KMRjo
n3E8jRgLT/WpAH5KnA3CjzHmYziBzh9O3epvtSc18treiOQumu1R6crs3NQ4inyy
Mju35Ww0RZ0VPJXA14yy2/W5P1RvxY+RGUckoqYxytT8+5e2hJMBz3jFru9jy5F7
AStI15xcyf32meJfSI2bfRIqPzIaRfmKtTzCoJ95gB9ljdG3C0WiHo4A6HMS4HpN
gtKEMAB8W12KugosCJjijVZWhI5PfHA1GcVzQaBA2hdUR6VGrYsTvl68NHCqCvfO
w0x5p0IBheZEpuuZIyGFyQQdUYvgm81i/YNpOYxzHIDUHO4ZDmWsLTN3PhF3XFjo
KA855+u1Q6yVMd25YZGJnwVXEwUJxmVhIxQ37BU54S3V8Zb+FPt7XluSIkVYmOyL
Oe9W1CqPC7FqKpLPzCNyE/FTKpqDogILcikNidNOWJlUHMx7rsiPAxvguvYsb7J5
wAylR7n+gCeUi4KMWWZM9T6rp5B/plxarK0SZpXkxUJInZkTGsYdRZ8WQ+8S6H1s
H547pxhmvNsz+M/+bBOhIM5J/M9M7I8iyw0obFNO7jvHC6xbmJilXYiyjcxevqhP
k9GCpgoQ4kdxZLaYrYftVWvh822l0/luRjNODpCacOhaHxL+dk6/h82LKP4UO3Z4
esaqjGU+6CUHb7/8cPJ/xK+nay7QQUg72EbVZ7CL1RigNGV8h2d+mgqSk3obZpVc
xTdCKJ35rAVscP29aQsgcF162fFZhgt9FY6SZ/9Tqr0Qc0t7tkVMq4JiRjc9HGjO
UXgEuBUoj2NNpeXrNm0agXfYOWWlWhlVAGUi68KfbkkrdERkjqSJDoskfBwYPQEi
3E7VTomc0Xfuo/1QXgRqSkDTlTHsXw5dl4/AJ3lOuizygaPxCyBGae82zcSirdS+
RMCcp5jyf1+600oa7njfqaueYnTOGA4zZmQr7gEEa7ShjLBipr5xHAIgrWEsQM3l
/4bBg0pjlSBiXpindBrbyDxUJ8gzkXnNAcyCl/XQr4Z0mB03OvEgNED60fBr/eGr
luhKcqt8hVzFevIDIOKYLJpODa16fvxUy4u9iPnAG+jeEIK2jkLSkFsX/cUM2hQs
EDPXBfIK+tb1IfotW8sfeYuCnzTx4665yETwgyAnPHe+I8Wvv166zdjy2Av0iObG
A5/2AELMk3CIYjvBxmd084Nr+9BIQ+v7a4BCMWIFbIhnRWtvuZxqO44Cyv7sJomX
B3Q663nbLDGyDaQbaOwi0PZ4HlwUx95k3q3krht64Zpe6nImRBrFnurAAmTJIsQs
kmo6vTQIs4aK2wizyQr7+3KUoqcl5WpLIiO8s73L+Re0F7PEJmfPUyOf6Gg0Zu00
Q8cANBk8EsmGZdjSZg8VRe9TolElyTNbAb6j0E94ClgiYvrJbcfhC+fcEZBCiPHe
dC+HRvc1leCGyZuCgdbYb12Z4M+W5ltmCbiXZr37yjkUGQVmll/XAPrhwYniiifq
1a+rtMwhSiAzTrXiTWexUVJ+nm/2NiDXnhBAxKEj7zb4JkXAgd8DFyYhkJGtB3nx
GpQQ+yXWAkkAXigjw4hFlnl14qnTj+ukVFUP25NwkzZ7sWso4Q/YTXKY5OUUGDsk
0w3929vY9xLgaeafeJVP6fV0eJprG/T7nngvkXsU34mkov0YuoWYvdN+ni7FCsF4
K0T0ka3eOLvl2+CsCsbQI6Lk1ZRsnpYhsTVy/A6rSiHMvBJxALjxXdMlD9vVJBmG
vNz3W3f4AcCzErD/fZaHJ6MtJIAyrqImnEjyS1Zcm7xtMLxdV2a0wW/UQURJPW2A
2ZhohMxa9meRlcYfbh4EKy8ZtztoaTv6sjelJD6/eiV6iR3cAoASidJ9o6LAgUv1
ophYjp1AJhwsSMnI6zX9C8LodtLMcvskM8UJKKt0fY0lQI32Idav67PfeUbmVPUO
0Owbs7MzUsP+cPHeexBsggr0sM2i50XfqO71cD35ayjTMBgyJXV8SrI2bjtipMmP
7Rzhhm6ybdWF5eIn6xBTyExXb7NEsFJyQLyLA8n61COCda2/OKyVoaqs4JWzRrOI
sh5pLldWwnC6L7W9NOdzSoHDXEHge4HZdSLeXcXHVEW0Ohp3Z7n3D9PUPwGmkCCB
59t4WvRv8L0upgOzusMJATqTFhgIejdqPlOLOcXEDgpTreHnpRdlLiLNVG1mQE+R
d4FszHd0BjGuzjRz7XfW3zifM1IuVkW2QOK21WI3WIf1AcVVFRSb6ZZS82tTXci2
9y+KggDTU5pk9Uph2npsiFihoeIDwVXxpJyhYk7wGhK3FHhSGlASnLTmA8TCPu+d
qZRICHM3Zdlzd8TGXMXZTpPerBn5Ct05hDl1UkHfhUhdFprgeiWq5VVkoOtuzdUg
BoWAmwzzW4xHj+wdkN13j2zykzU34g2q/gFt4MKkyOpQiOYs9HRQ3++pK/hrpWzR
yXE1ZaDVuFSGquXmJ3bhVwJfGhivxL9RgmYKIzwxONQNlNMDTcej5mZb2R0XO43y
CIFv7HvXdomgnAhbI+ewbV0TqvWgae2S2DOkFZe+FSO7pwR5qe2rHgQBq6kueZEI
XmtwVMuaKipYLD0IgbTjGQRjEMVGNWdSPtIxUZgNycHw59L0btfSG7OjgVeCVkj0
7/vN3EY/HNpmJERPtDep2371SBPIpEFmnaLCIophiiN53/tBOeJRUOxpcTXlxCKa
ApZf9h1n8W5vjyrQ89HPVj1DzIik9A+6seCXkJZCzcA/rvdF5OrtXDSOo7S9u0xg
rToOUWwWS1Wat3qxRFXhiwrzmf6AjwvTSccXvcRRNcidrXaYRYBRfnw0Ltd4vgjY
/y/rNvHf/0srIm64oitQ8Elj5O3SffQadk1m8S+LdlCAQAsdeor+V6+RvhYvezxj
dADyeqZ5i+yLAcAmYDhvuuNBlS9SBzNZlLXtxVNCTtVQY5ZmSrKvWatWcSZkbnCB
ESi+Uo8frYtqFo8vXlQf+xVXCjAjO/cAEHEjF9F6Cv2BYjJ0HA0V5purU8uIjvz+
UR4r830tamZvWKc5d4tRkMhPBPNNXsQC5WiWeCVNvWBj5nDHqtJIwq8vHoh7gc36
yISCxHDQ2duCXk1G31amUHp+DltE0HVpN2P8cQR89eaNVSyMMNZJpnHBnDK+gT4j
TDIFapnbF6yW4V0A+hU3Q1ytKgCbQlp8wdjauoQgLPJ5aFNUoh8TlccWFk/kYYiG
mAoYsHtP6kouTSYrCtodlVBZ/sLmMa5wPODn9FUOMCaNRy9M94+DC5SjMnbBaCEF
UkgsmynqqqiuzIV6wrP2MXEGUP0bdCUS98XzzVXN1nxC+cUehYq8qIHb8yVhyxjH
JHx1ryZwJEiiheXBdSlYREXj4iQ3poYFe2J5g7GEbyqDdTdXV+O/bPI+6OgsXoQV
lIlqvl2qDHASzGaWRgurrlpSjzzOV3xywuBba22oPJui5U1esJXSyVod0dcQQo0B
6gw7CL6nhXRdAFc81hSOtpnpuayJsfnVRj/mqKSRf9DdIZxQuYgYJrKnK09cY6IW
OLFljhGLXHUh4fvAQZHp9aiPuMBmcyrNWiiRnnc8hDsrhOaPKub9PkstwHC//zPe
5NcUw3l8Y92AxzfGGu3NhYVYopS+1PxCxc/YTw/Ay7myc5AHjQq1V3R4qo/UdwjZ
jaKmid39JZ8pmu1SFaWfQFiwb+q+QPwvJJR166QXag4EEkfAsUUWJawuJbzlCyUc
5zmAeiyBOSiBYTK7gYvdBeoUNMOfyqWci6vsrtBhvw3cyg0azV6kkSVmA2z3MTLj
Rwcq5ilMO7A1g9qt6a11rFUzV2v/vLA4WOX4RDI3Qg+dRpZx7F4DgCNMGr2LrchI
zMOPdO+Zv/e1YnTDnkmggepaaqc/i6eoZ4irRVWRwSjAexkytNWvzP3d6pZFjkfS
PpkqiGBEs1qoUyGWhhvJS8zrQYYofnOytg0eSHZUy2gGs6xZhfIEbz6FS6hXHDmI
hTD3UjCXexWS+EQ0Sdqf0axwvA//7CrcyoCqvqMzqhzfy8Hn4JQ+S4Xd3zP8XfAl
4+HIej+eF3DZyIqWDqzO3REzbWCQVRbnKBMo8rN9H1BT3WL9rpIN+KHxZ14ozpol
dVs9oDp3M7DjRDOWMAa+nIe1Zt8l8h+7rZdehBwXv52OboMU4lnDfw0fTa65ImGB
q0b8aOt2MBbdI+F9Y3TcWQN8UAob+8F/JdVRunL59AV/SbfcB9DH9bzaoseBedZU
Fc+dEHVp/Q6BnKXCESm1U1oA4bYaQhHgajnlLsyD9nlubIoepgCXtctLJdsBIKLZ
P6Fak5vrziNiqeC84KC/pNLFJT1Y2ONMubAzlS39gKEtuIoN0pk+mNSTd4UjPP4N
7ROBCIJRPsZ40pyF1H7zNxPh3Uioyo+88VcTzUM3eqviCpSeoqtH75FiKJ1VcaFs
gMwiszavE97otO8/s18IxWfSxk+619WXBE0PWlQ68aHEmebk+UdAbG9sK2Ul7TcR
OwD18Ynpq9FFJPgSr0IIlVux+QEwOiFYjF9r0EWDRvFxsQUr3SOzngQJHc5URba+
MSMM5rLQnOJeU9zCbQvJbfzhBC1Ld7uHB9uwiLCPY23ZnAOtfx2Stg9DRzF9Jeh9
rijJQHfqLQCJrFJv903XMz4hHppUTAa+rWyMvoMaPWAQBy0DhPAloeD8y/dm92aH
J8MYNR0ENdK4XlbCfnZn4LykpD6O27JOhVB3mvkqqBV9j1gDbjIhTR8th4/x3TQj
2KpI54BRroST2BuiuYCkQt0Gxef/o1bqlO+TE3qzD3eXTxFKUV95NTTsqmBugMa6
VRxpgG37sf5npFYudt3YMwtA7puWFXL9rgLCXlus1Ws9z3sS+8uck1zQ/TVFUOIy
XmXobzElIlM5qwxRDk9T8UlkJJmYtoAo2SvVXBf/xwZBHLJoOD4Lo6t3Ax4/tbMP
KnxBcYRH8+NvMmtvnko8J1XG74QZlC1laeWu8/49GIQ7IMKvJaNb7wxXONW8c7tA
Hf0ou3jnNaIG8MiU3FUxD2QPTwvl0ECX9H0QH+8+amRJ/XLfiU/mx1SUUJIEnOhh
m63LrEAE/oMHuztC93QhTUglgEjyJdc1QjdWJy2GwUp1rmFp3jJXvbkBCDoJe/Fz
+pUC2Kr+RMea4KJwl3kizFJF3iCyiCga7pfGeUTOAoT7fJXHLi6lq3nFBF+Li5xr
fWzW61wzge8hNK1RXjWRFYi9DDnFE+VnZXs9Opl44Y1xGXwpDm2JSw7gNgRlCyM+
whBhRi2aJ6LWVZJIvk5+FkXId8ndJCW96hXCyNOiLpuOg5AoAT3+3zJMTVa1kSR8
QR1USO7wiOKCs/G9pZiSfEt8sBOsLp4E2gHz4iYoZRMhCSsiRbbGKmvV8d0KdBcz
gk7hq/VesoAro4RzBr6K5/oSzyVL792CxmuvFuMC32HPe2Gl4BrMW6hA7Znn7qAL
ZY5FzJBPPIzqvKiBh6i7lVmrH1V+GA0tJInHoAy8xGC5f+yEXQmDu/waukADioRx
WZXRDzXaQIyz2PLq3NelLWSVEWaFdPaJ9AZUa1vehtC0yzTea7ibNdypMTnfXnmX
AZHKnQcpGiFQQaWWvx1Lh/gRZoSKK+5J/vqXuS8NQ7BmBXwmHESHhTPBFo4S6Gad
dEywLRotKojtaAGi5JdJbVgdhQMFODs+JviLz9/3CAXjDxG2i8hsfgSeqVVaRMGp
3FWWv5yfSqc183ZT8VfCleQiPOVeBvjfps5LjdxpJpS6I3SleeMmCf+Vp12ytP72
ij39wZpMCxuQlyO7TpYXJedZ5WSEOCuAp5I5hZWsRs5OTNoOPTddNfXDAwNAVu6D
xMMTkopOyLBhplSbbJD+EDU0hS870Pc5UYMyAOO4M2//qjfWduh1MtF5Qi64sQaa
0eKiBu4AJ/LjOpRrMuFygB0ZwF6vqpouiU9tTV/qodl9bCiMdk0jCZyM7mi/wX9y
sFDCFuKYfTkCa0RprsFV2CuaN87+rbxus9dGtWk0zusn0Ds+4S4YyhCL3BBVzXrz
MwyMqjQE05RIb+M/ebG5lW4wToRCu1++xZTQMcCDvYuebIr4M1/ku+5dP6+xzMtq
hb/YTLHB36CmDRWR1pj83husC8wZL+PKYiFmm46tpWgkfEuif9r+AeYGbc2raqNJ
4oKoiSrVg2knzIT1GLApwAElZ5UaV/pHvb/lkmsw+OXcQQHMWeYYWfdk/q8gd+O2
uJPPOt/7xvO8XpZhpcCevhLdguoeh4O5fyRoHuiGr6GaMb5iFlYdyahtmduNWXDR
rtMBRa7M1Gv9ymuKe7FrohGWViPkI2OE5FrD4N4kwGSyd15CJL0bYET5390Z/rXQ
2jBuT8kZONq+frN2H4MpwY27KAjTbXdp9WBESHQhkgsFzq+oV77XQoMtTw8K8lBN
X29+aRcXf6koEYFQ15lUnwMlk+dFQ2HLb5Kz8OmUsFYBdVVrN+to3Dwhx2irco8G
qzU0zfacOk4x3c884tvNfbjPJ8uDCIzGVq5MasP/B5vvdVLrHD0BnLrF1tfeRP3h
Q6IioGFJdw7Mb8O+X0mmFsRgcvTa1/iGvAQKg6aNvjpA7HwZS0heczJK5ipGm5a/
H3pHJjI+4oG+prhswkLpgY2uQMfLcI6I+mxiYzp9impN5vIsQkIUQWPcBmyeHU8a
tIMzmBdUT2sSKAsH8PmjRUYmdwIxJilWzNeq3xejqo0M8GweMf/5dw8hImUADen1
1F7h2+oyCdLh6DC1s97gjeOfxcyqKvA89Gl/BuQxeLT9IA24kMoBgI8n/LnHZ56S
1P7FRodDQeeojKDhBDFY4ISLWNt6itiU0xNjoUmn/zQroC5LCnSkVs4Pj7jQtYZa
xdGcMu5rQcLxCAVGpmFelalQy+troHtpuQfx+DX0ebmnMO3GeBNks2WL0CGty8Fy
0udYjTx/CWItqyeZEZT628awmuNoVmtOzXFw85UysgtuT1DbSD+jBjO3SjN5r8w/
ur5Cj4occ2jDErsIzFwFFltXWKnNvPPy85iRifYY+Klo2WmC+rt5bypo4e0NLJ5M
F8NymH7awbzrmTzUlPAR1htJ83UlG4DfmRngzth94iyarhiJILzzgi8MD/iGJAn4
7s1CqcC1nPZnM0fw9xBdo/0gN4SP8VFHC5J8+LCDrPatLk5DGG7NkN3iXKM0iaOZ
Ooj/ukZhEmWurH+5yczA9tuYpkpL5o/GmCpN8RuHKAiRim7IjlWtWArWfqLGrIHi
ZLXXoNo+7XTqDZYE7LRn1nNfYvgSKdTaMV+DSTmRXf1lyx/pqJ9woyB5W0RvXK08
D10h6w8yno5vJDq3YfqA2MGQwo46cu+mWLzsbsCcN7EIJ1Hs4P+N41PLIyv1vdCP
CRrK2QylITExi0XdD58C85fdAYGMacla+8hex+f5prOrRpMeqoNAFiHu864An5+s
hcl6XZyWZhA5AhdMcHmcZ1a1tP44BynfNroHSl6GMQHoegeHP1izG8aw3sogHJth
DjGLOMYzPkZUvOzTCHcHJ0Nf/F3c/37FEyOp9Y9eJBOKaXj2V3Ful6bApswUHgEx
JBeegWO8Q5KIUMbpRCWSYYnAbKq0opIlcb/e+dChBwlIGqa9jHlu5PRT2tmrSgiV
GRQWidklyLL6GtuLvHXFl/QdgAoseETy6oxyZXIRNkZ3JewDF0W/+x30U69pDMaa
vsAcAi839O/H5jE0CGECJGvLNpLXGJJa19HAUm+Akzln0RJd7wugAjGMY8uCJu6z
iTh7iZmcwSKthhqYqyV9S/dlxaJ14DShyhJqFI/n0hkrFrcLYkNXud8rRYk99dP5
qVeh7zsOYWKDYPyfnPbd2r2qocl0KSU/l1Tu7GQy+u/ZzCnhsXJckQTUKHCWG98N
3F3DKSkbW1Dxh4RqhG2SNaBuquC/N+yqZiMreiuzi6cEDUmMOqFdb5mnvJDfpEeN
fK1K/2wLoemBor514hvMTw0F4KP4k709ZtDaTziyswt8s2B8Gp2JybxNZC4dSTiv
d4CtcRlPQY0vDSIkUe4cfyg4mBdviMU+nUORYRwfQgXXpXt/ptH/ta6FZdZE49Ia
2m5n3qBNkn8T0Bpo2MLCNfPr6SyS1rZ9A3gMi2ZB4ctYgc8kpWjj+DoCa9b7YMqX
cABytB20j109oUfNTA3UluMP2kMuZzAjaGR0KP7NHUdwR1XdvaOP5vXZ6d9k/jDs
J3wVx4pE9jY+T8hvJSACX3IrqfxLzORCLkNneDIqK1UTmSgE57uZQeF6dl8PIJFe
ywKr//3YePrHUaok1k9awwAzgGUS3oUVt1I8x+6zf5MiryUCMSc2T4wzIHmjszc4
ldjKiZvibBTtcF3Qu/L5dRiK4yqCxfKsLBkHKxMPNM4hlQiN0n6PqFih2ZPDulVl
jZ6HiUik9+KTil8M0TmKaadjW5LrX/BjYFhOn51Tm9VgW+ejZw7oELdQGyeDYHaf
5vBbPvBPIQTad9f4o2veu1gzjpYJzjqNEmxQFvGWgg4BbWH3H5TUL+xL3u6m/V6V
vRI0bG51IMhE7p9SQtILtX6ikBF/UXJZhkRWyDQWO5/MKqL/vaoP6KfjRCRhe6La
SNH9S2hrvDTWQWWg02tdYIHUSz6NFSNd9G3AMgNr6n/DLFBCFAPXrbYP5+1KGwfc
ESB4zZKlmTSYdHjTD4tcJaWQ6R6aTOVbD+X9JRn49blbAYxeF0ijuAMVjaum3koj
e7fHNeNMTOGBILwl6XzN98Wb2C9wBd69YZqTPpYkKnZiH4roCYowXviOp99geIOr
wPutwENhVt98otbp7tAMXExNNHFljGQCw30LxyozK3mXbI8y1fXj1eyBaxkU+jVI
lv6VYtW74bj32JHyACa4BmCaqtSse54KyVZD1nguWOCIlRyCB7iYZWvJAIGYrBij
2LbmhNCNx5A2ejta1+XGhnFiuNtBwlWeyOM1Fnpokh2DkXekMw9w932+8o2RqEd7
L6WVS2YTSb5fTzp8WgWvtHR+RfS2QuCibbc26F+JjpZyuZz7AMTHpU75gr66Qrqw
rGEFr66lNlBMsrr3o2z4xQI9Jw4OhQ3aHiQ6tfeTWUltU60H2axNGR+TjgTfD/f9
iYKFDKK9Q8zzs9ilIc4BTaqskBEq/Z6n8J3mxMppU2nJNOkk++2Pvb4FKo60leyd
H6+EmFfTch/7+LAzuRGhMvFLT8ufrUYlmHm0+cIq7oC6sEbtj81+EHwh31tzrXkG
ftA9AGibAWyMCLnhDMmIHmIXP7npKit0UPDi15i21SqWrYB91epfQtsymrn6crlY
qk6nYNxeEvZVU3eSzAPiDqm73RFrH2PKGjxLJapHuouKGN0uuQRgzVQK6kTw2EU1
DeIJni/RJcY9CeXsCda7pZo3vmkgFmLFrGviaFw4IdRwgbf7+rrFjnl/gtxHjrHG
3OB62Rqa3JddfyWEhL3EHDYCD2B8WUZaVIiOOILGAyFDmS13SWw3ozGZ/Q7GEmWt
Y142YeGZdMpXWtre/x4/nT2STJqJJRMWZURywN+C2bGv5gr55WZw6sDJxgR4c1DR
GH6unjMlMz4HirRJi9GXi5c3AmOP3FFZwzjFf5nf75DgTIlDm0h2gH6LAOdLMBzo
3LCb0GFqcmm3FSWDuS12cwA2A0ebhKdkGwuUidtarHPShpc+n19w+u8Aa/EzwlOP
UNCG/fUCREnneYNJ5J6ujM1kyxTJG+ZezOgac/SOdISri0f0+ChAbg/7OJCpzHjM
bOSqoEX3mOTYz8Uo7B0MkZgas9BJqiq/MG/b4NMKCSU32gYDhihIFwgVINcnMRyU
2t9VIBZFLS/bspQnqiX4cC3BUMJqfaRk5n2eaVL9KmR7nTOdIUwUYzGTMwzmJAHn
/LS5h6Tr9GH0e0lTuLe4Y8m9XCMTDiKfjsz6/05KW+BsGsrc7018AUD0uOb4lXoY
NapQeAwoPtlRxdWPBHejlmdwOqhso4TsWnZh2JCOYhjfaSuoo1mlDmty0wQl9n+B
2DHzgCNTkqUpvtZ948nDYTHrkzAQLvVq8Wp16ZwEN8lTOAdJNGFSicGLIGA9bE7u
9JHxygDMaYn2f8ebREZmu6MzO3suVuJOITE9jK97DkvIaznee2d2g2pX8fQDSW7r
Ynk4x1YNr+lP0IWpgLIx+kZdvYzL5+X53Pq8xa9f8S/dxDvj9GeB5dCWx0tTTx6v
UL7EhwmQtZGJAUBLDXWtudJ6zDWx6r9Ie37LbDjqQddAwNRyDBzAZpeglRr22R76
yg7L6sviO3MyRekv/f+BZOU4uungznrFfrY/PAohBn/mOUJSZZxerEOwUVQiHhD4
wJxVKZ+ObWQaxxkNvzQxA9evuxVJOw5EfX2uVv1rxVCiPrXnX2Bv2nZbAeO7F8xH
nhfT9a3/4qjh95PXoF6v6eSALuquJw0h4Y1yxKQ/CO2Dn8wSMcAh9OQ967oWERge
mx7kmQpdsxVz90ZesSy4P7xbNaOC5sOr+rJW9RhLBATwBJzANs1vBVvHPlzuQgO0
c6ZMd1NACY10cd1Th6q7PeSlBdoftPESIVoOtD1kQt477tZWQn/i+KKVXwdEhxH4
DTnT5CfeE2eN0c85Vf6//KU60paaV8eOmbvyI9BjMpdSXUYDYGAkOe5cht8f6qv+
hKOkuPLSXcDsi/rTkKuQwXp6rgmFpF4Pgikd1is0ae8PeLIfAUtpNSodPFpMnw7l
ky4VBQM05G5hucb4rqKMGZTj1jkgzoj4eW2QyhX6mgnotx55MMO5P4ebd11+hp+s
3AE4HaX8pXGS1563vjGrg0Uw75u7wumxWd8i5SVkE0XhZ6/MlEniK4ABXb2yBX39
tAlBeNh72MO4G6H1IFpRcPs+Nzwe21YV29724Hk4a9TWFunw41nD44CiTpZlqHGP
Tdtu2ECetdMxIWrTljIbkfJVG5Za+uAGk30lCLVMRx+TYLoA44AmAYp0WPuUZ+WC
i+X8VrC5XG3QNpYKGQ5d/alSpbor+Ch5scaFPBiZA8Byaoj6qHlnK1E1ERaSLpiN
Nvur0lb6VHYZmCvS+jHrAaEFJWbysu3xoKI2INeEmk6TxU2bZXzNSKek5tPGNFwV
+CWv9FvBIvD94z3CnmVffFixhb7svWDDv/GFydMDRMw8zrc3xCEiM+QkYesUFFvQ
oviJtE3HTIjJTiim+/oBqliB/Yue2LsvkVnRzaJxv7ycYIVMdJn0W+pLddbIIxID
miXiG++2hWOLshoyVXaLdj/2m7TIaikpikIOqRkyzVsz9KpwIRi/02HJN4Y2Lnch
qjvnCPHr1Xo7NYJb3h+cSAqL6fsU/mkaMcvf5dMgXKEC7mqgJqGyd+GGcg3gAA6b
ZPjYATGmTQ53nLhDKFHYJi+5J0ZVNkgvALK1pKbIEjzTLBuPccwEDLoNwV3qFL54
+6v4n8UW1eDoP4cOLJdfP5jmnIBim+4ZLLXokJrNkrAj3DLx/XN46vvaWJWU3mWn
l/Spaadq5GCp+N3GpimLPMrGl+MNgaq4aGyPRVKc7412LAuCIp7JGTRGDDbg7JUS
EwITKTjmqiHkaqg64PP4wI1vQa8zDfY6MfVHbBZkxoJZR+IhNdKpGv0Bfz2d1fZi
U8kAHYo32FiYdLFDkKMPz53OVV7I26bHsSd2vW9oWjspfQhAT42t4hM6iWcuZL93
CmkfWn3+gPia44rtUiEJp2QDqdlSs5AOJLVCZ3L7myLdZnrvyHqs8tg3Rlyys8cZ
34dw/uHgCzwee74egts9WYGKMjy/1B5YsCAj4jcuIJMbTIHNl3x+f5fdO7+ujtgV
2jGS3OvV0f2aF42TDmbmI9f5IFSBswFrUD2Dheb62vLV90etwlVQZzl+JaWQdvgl
S/cCqn02Qcwa8zse94meyTrY+PLkrlkUaeXooNbvGnLVmJ0Pl5bDuIMMTOPzALw+
yGkln4F0tT85XVS+P8T3XEM+1uGlWAJeGTbVwY1Dr7DBRcylB8tHoBPT0cSZUXwj
r4icQ8F4tkvGMQD0tH31Nm6SCL3c70e3sBf47otXRPT5PiE1nUKzkMzu4Rdix/5C
XkQ0S48gcsOTTr9I7hefOR8zNM57zlwADjrR2dow1x80ta4/dD9bo27OBLeUQdJc
M1AxOEx5PD51iIT/H39Gyud4avpPTTQn+rL+QRQWIoUWJGtej9+yLjafikshDfFY
aaw3nP3AWMJ8TK3gU3DQUwBJtnlT+TeyFtql9R1XL+CORP8+sWieVqYwNstzuc0U
73uFLbXyOoVTrma3tJR1K5v1BFqhuxuG3kqOn6iSgfWpDEO8XHiscJeAPodlNffX
aDv02+a7/6ZmxY6eaPsxMkeYuCDj5CzWEGL63yntSnXKAmWPlzmDMT78OlwnOiFk
/evl+aLpe5kRDlLt1h4Qnzzs7imxkIERLDMrbe2pYuo5A8cW9w9o1tYgesPc7mPo
sYa7c8akO6Sx32K1eyfAF+2JCkU2loVjMU0SxA8VhLZS4/IE65OIWojkwCB/xztI
HsezoC/lanyRVIafKf31qTiob2J7q6/ZKUcF8Ai5JXdDZZ+5ajuVU7/ha4XSRhib
MMCGjd+EdgP1/mFwVEC5W0aoTLFrEGeF1e+5eN8REnbQXr3e2jEy0MtOcEZwD5st
+WazCL0UX5QvB98xTC8NLQLJDAZLZVFFUUEtJa3ujC7fgqMZYHvHZ44u/T7mGgZY
bUxot85aTXRJ8CspKxQJWcOmHVROfPc5uvKwhGGBxcHtfF/A8RwKWZ38nA046TxP
fNRU3hJl+L+lcfzlUzt0bUpqVLrw6ZTi+UHWf8RNL+WnE7W+RO7MdL5FS/NUjvRO
fhqxWyPgq9hGXZ/fL5VvAXoJklpUOOGRmWr6nks+OXkqOhQEiiaXjiwVdW1IlO19
P4s0QuYyaaSRbRsX8tDZnaBk8W+dcjRzXZmzCtOYpElch7gkumfsg2Dm6WYqnQmZ
+10IubOkIncENXtlrmvSeWByxzzQi+EPYPEzA0qKDZkK88de0qBf3kvEgO6zFC04
JoXdMTPvrbny8nKqvEfiMfkGr9Uf7PUFUPWf6meLkJVPPmUr0RrZTkfwMID6xAA7
3XG3yUPJulk/LRknWiWYBRH0mjEy+5Zr47+S5advrFY7QIpLEwmwbYoSbxD6eeJh
KWsg+mwSEGZqQ/HJCF3j8Kjnl61z6VpiQgnEigTFiIg91rrFuH2YGAn/W6y08721
Gdlx5hy7T799YsH9QFUWbboT6qNxALo2IvLsCqBcapgjvt0tFrcyBURiYvncqQi5
hz4uJllNB1292cB1+KwH7j8y2pXRvGA2liNFD8suYGO8b2A+dsLb9jTzIlIX3vJg
b1mfiPK53v2LL/dG1tt5+/OT8C86Z7JqcYmo6yikqpsnIWqIRUmteU1SXTbVlrbe
11HHs7o9gnRyeCnWQR/X1dPd/YFNKflVLWRq0QnhA/qrUWNLywg86ecCc+AyNSTQ
KT1FkrZ/kn8ac7jxkdvVKSj5hBXv5zlExx6TMNoF4NCL2Aqfd8q3ip8i0ld7vAAP
8drEWdcPpP0MIJZIpMZQcZQkYvU6ChCuHzJQKDReCT3qfaoieMXvh/iyJizORx6j
ipr3QQ79GBIaPyQ4Jw/YDgEiYXNa88MS9skaViHvWbZCYPRGiQd4oZDSCvTD8lOB
N84n8A0WH5NW8gcsjbPmX4Izk0C1btp8NjB5RSuTT2J/LLLqgOQuonGyEgicttlL
2V3irR4tCK2h1UVNdf2IkqguKZi5rtfI0WpuI/1hOWlKzfY0hNrdJSe/f5FZiPkt
woY6O0brsMPfkNW05pOpHs+m6IyM4s1xOtKcSIfy6OJX5/SRXC5XpD9O25cNV869
3h4g+e67o1AW7LwQTQobT98fzG5S9LUwnUTDZldkkNaEl+9MvRpcPPzMDkaZPvvy
mzqWjXB1eL9w7TalhY3DS9yqqlwNCYA9UoaPEQzFAFmet4SFYnLc6NsVuuJRzHHF
ks/YdTFX3AUnJiKio4o78l15fo+mdbyZQm5aIY5yxsBtyBJ7O/4XpLOU5PoD8jYu
cIkXnvopn0KvOQNSWBTm0aSQPMnCQliLmrduTSloBq2cD9tUqRTOOHqnlVw29V1G
BuBq3uVRE8m98SeHyTOpeWPPqo46QQqbDdSx/WkUlz2qatpNo1dugd7QLKjjZ/6r
Yv7/clueplFA98YcRFsx3dnoKByHbNErjOz2VS1FSQ2av1ZMlfG7u0v/tZfMGwy7
BzeZzgK8rnqhf8UZ7QtJL+Tsb8SdTTZqtldCxA0zTh3A3mOoLP11tLECV3NnbJhI
MTESF6ZotbbtZUT/csQsGBtUJFIrJPthXdNKFkjN2rQ6HQWEnT9tfyc5/+Bm6az5
mhm4tdT9od+3/i7MOZN8j3eG0Vmio9nTcnMmfzXrBSobbQtHBYuNouKaLAJ2gEvc
aevI8t4YgAO4WJTFY2HW9Ossguzm2Il/grvfhVKeVwTSY64aFnwDh3TOO7k3KApY
pxdrM9fUvcJ7yLwFzREV/V/K4rgTS9L4DPtFp6XX7yRF8SQ9trI4r6HHbe/oHPgB
55pXotFZu9npQXiAkwgz6LkUy+ZU06OjjsacUDKiRadP3soLKCQMM8dQBq3B0c+v
kdGjUcdKRuPU+vQvpQ1mwkMwGg2PgPoAzUzcZ+NE7a9uUVM8RqlK6EZVa9xMzufO
p4M/Is2eDXUOXr5YlFnsWTrQ+bQpOmta7Nd2omdfMEr/K9wDG6OvRRZMmJYtY6bU
N4i9tv7NXUZzzDpt942zvR5jixFASbpcLqhtnMPqRzK4yKkv+Md9Phn9QI1prbYf
NOY11uc7XlDVMB6IGg07Vlx26ZeCle42KL2hvLmzdPLZvo4Xozod5v2tJxxBiqow
j7S2h2fyVHa+hlqoN+3/TwzEXTMakEAXGn7ymESFGgKh0EqXiiPAdmHhGPVCoaqN
h+541jbE9Sp1y7zSUXFrV3kKDYbZTtCkIO4cYROBp18AoOahZCg4/bYZKNPaqLrb
ftCUHxwIq8m3mdT3fQFI+LdJiu0U0YiLLpLivLE3l2ZZsP+10dul3OOQ+BDsfD4h
P8pFXztTCRidCkaFu+bdIM4zs4wB/MSeoyrcyktWU0odmVk87z2LLQt3bxT/plF7
ApvYT14at/S9W8r2k5DnsaprLtwXqQUJKWjoffc+qwkSgEojR06sofacnvwF/h0A
qxdXmEu4H7cpxMLSUuoo/2HkqfT71UqHEu/l5T0ZA0hOPUIu3jufye/DyDwyfl+v
0drq4UhlE+mzvOdVVVYHL6zZYBOgmT8zLxth5MM3aH7XngEYQFmIcQB1E7XVSnFi
wOyX9zdmeDGOKCxNyZBMpzN+kNLFjSwXCS2+DJMUNGY9lnpvBPlzMImbFho0KQLd
/TweUmOPRcOPAT0iEceSBkFXq2LyBwC1FUO3JaiP5i+Xsq2Tteo9THBkekc1lBEH
71CLhyIKxJSUVt2ZcjfFWdoKQAPeSTPJjKt44yPOLAVOfFNQG1amhvk8CT8YldPM
e6JnPyFJwxCkpeJRE8/r+ecRgMfV0J+EiiCaFlgM3Cb0+TOqsaBQJMGjn9G7PaP9
ctPg8kO8qpPFtaT8NdcDEsVxBdnLCBvftUWp5rPhjZq8pkLjP4mkVc2FUgMuTBfh
av65+XXh+8G7EQT6QQwq+7orpb+sK3DKGFb+WbiPbYYKgF47cYBgTLRyv6d7vssz
67CN+o1QxV3f2UMy9nkYOnNCMcuDoj/FkBMw8OV14XMIjtFNIZ5mFg1hpQsGtfqA
9AY1aAIi5WD+NJmfRMpmUoAwFCcsQXLFYvnt/x/WNhc1G8Ohyftk/2OCKs0oAERb
y0EWcuhlLJUiguZFogcWL07G0w06ri6XgcclRmmhoq3rKEoD6oK2jvs9g4c5j5D1
ewLTn/5xvaDk/fb+5uefcgdLk1GRA83N8aIb+OZ2/D52nvCPdHkKe5wEeHammdOV
1AhP32nKuzQbx1+PcuA5HcPgRWEb7dd104e6+7MfZ2b7XBWNx106ZvqTBecI1CCE
Qp2lD4zg1tAdXJgEF8BWOxZKvRCI1I+oHrVGltu4zjRVJnxWPNe26V5LPz6WJtJ7
Th6bdMJ9mZSLWclWbJXbk0TouZKtj5KOb1kNySCPdv3x5IILQFqHgS5LDu0dYv4c
KptSXwoQQ4FVZ0hVSGiR3cgw1ZtMM1Mpvm4r8/wxOLDVFZCsBGxF63dINCHrX+Y8
kVBfu0BzzefDejHAIvM3gjU5gJswcpcG3zaw46ZikbOWnk92xk9CCTAj8jv0tarT
3qLtY4U4GUltKh90QJXzyV0Tga/G5e1JhviYr82P0hl2TXqB3s8jjpA3vLn2IiJJ
JOGt5BzNxGGNa6FxpPuD2qZMSwt7kJazPQyBJIRH4X6jc+ycMSrFzQQmacXH0Cq5
cKzVoA3M1AfgX5W+j4BA9b73R/9pHACjozjULKAzo2ys07AXBGZMOL5RlNh0aa37
/AhAp0710kksj5U5Jy4T6LMO30waQFwUmEl2dOzHMahrdsdkbvWSJ/YIIeBFtHuw
cw7e89PUY5dy4FzkdOvA2uAtgvKjN+19GvbC0dpqHz+JpN9rfX322oPpFtgJp0yc
Sv/pX5JtxMJezG0M8WZ1NNvEi045NJWK1VmZd69e5IQ0DQXqHcOOPFQB2SWW+ava
ZRac3I4sN2zLdhdU7KJ9qI6uyBOUNrToDNu2RXZNMo11mvlPRpXTfhcf28pggre4
lI3YEinnbCLiNBGQ54045Rg28edbNcEka0rZDP1k8zW7GNMdtFPuZ/U6h9jMJbwy
IsPCl0Zqyi8pfmamFVXUi3E2N3H9xWjZd768HSGct1fk7msixKaAYWrzuVgTG1/P
JbRSucS6MN/1AqpuzVdIzwpSc3p21TZwUNxAIOSL1pZgpDeZGaoBvYs8wtSceOPe
B2NBGJ/eerIXo1UoxKVn7oRy/LnTKCBMVsnKy6E1+Lf5JLr4CeVyTr0AEzapnEfY
xOv44e1Uu3MhFMPk0/Kd0obj26zePTlpWB/Z7SEC0fscAhMjitxS9uHrObT1YPHL
1UsT1teLW1Sa5QQvFZhnw9H6czeY5OMtVB3GOHXicdj75yo0c5hk/qUTtkpY/baC
qDcoClw12Xn/GrlvhyKlWYdwrzPd7r3DuvWyaI3Rc7MZjls2gWPXU/SdlJ2t3rKk
aSzV5Rjjaz82CswcQOYvYkW+Ba6K1OeloZumysE16tmFL8lfJZWwNejUJEqiKOwy
F4fxPXtgDVhZzA7f4mAvzv+ar2oY+v4OKJcnrKfH5KWQWtS6/HjVK/mr8rEINsPe
hX8Ilk8b8qtKFnsUf3aUZyf/TaKKf+LqoLododAwI+ktw+HYqJpyRiG07ibtjVpO
3Yrhd3EIJBNfz13RmHE8TB6MfKdvajaZIaTzE1J6fSpPukSJos12Jgty2YTkQSOq
IGJo3O+Wg/+2+urZ0vByD3BHcnHvPVzStEegPgyFczLLM3f5+IDsdCLTIOUFI0+q
vYnLDiX0hDBlq056saf5x3Ioza84M/D1FiXd34V5GaslsKynBZYk1CJoYTkfTKcd
bd6O62w9fAYyqZsa0aj2kEr/pK9lnfljfGUa9K4U6LcsRbpEEWjy09I47i7jiBnr
onBNZytc7GzTtW0u1klyKsbOA2bvFtUsU0X59sC8nWWUkldtlR5D0bx7ZQnBRSOo
fj7MDPrySi6+EPvaQ+ki3mVVum5iEUBb2gObbWbw1+Ipo16+981Ns+5AeUCFbhdt
a1NfYglWX/JX/PsGQ0UBhkqWuRu3HPnsFLIJim+PrADbcCNKQjvNAhabq79hrjMm
kA926849upp/pEnmmjYxHIX7BWu7NLmaLTT4kX8/9+yYnxlb32hT1UN5IN6dAIZE
zQtmxAjZqk/DVOwyZDQ8cRyetiMDYWvdIAXiLRBFHvObC2WrikIpNiBeljToKkaT
5PQtVfowDqZU0es2Kcl+sxAVF0C+RCHjNSXoTYq07UZliwndDXISzUvYtYetYh9g
gS3fGhU12eq8Hqw/pj3y5hE8yjlWdwECyqj4WhtEDgOxkBRxRUMVc5kYwT+omXrW
1e2KAm6lzZAWA+yo1mcCspx5SZf9zmjFT1TPPWhbMIJhDBCmpraCgxOdmNV09YSK
on5F+yJV8m41lGVEpLhOoaXvOXOdjljHH4+E7WIVfHkaHsI0UUAuI2GQgmJOfTPm
Bqg/+aao3nMWzaHq5sznjwSeObKs3UYSEX/SVLULDpVSg1T4YWZ+zbpdgbrRpq/f
iGC+YoddWfxZVjSeAntpgbAGgxEwGbjlehigwo+dBncNIimcyuGh4piCixSOvHAC
7DUgxqzxVnFBDXFFkRiNg4W8xlAfQDV0fdmfF9p42DbbtbdtKtWt5AA1kooCz7Kk
pEmvUVtlwCjwe8fXAkza/ZW50yHKglR61f/UZv4AlQR0wBI7Rm8jWtQQB5QktP2K
evxCrvhCh/ezrSgQXjHu0awr9s30p8ISd2n8u428Cx+scpB2BFFsNaoTTlR3groP
GrwIQr6nkh2U1N3IrM1TKajzFIlmJVUHJ7Z58eI5Hr7vijNGNHp1VmVGRVhncoIN
Bec5D2oRnoaE/Yxbug6Lfc41t374W2vM5KMT1sJAMPm3PBdFYuQZCsBiz8UUmFOl
qXq8SI9GD31F542ppyjF97GZgUcFMQ8SYvkaNNOdQms+9DVQIZLsC1KO7rv8Jfda
2roCKRwISVeR4yTjIwBWiMXAbB4O+N8018Ge7aF4QDchAJljIkXK6+XFObvwIpki
4tr/PWXdcXZcWJMpcTF4dmNjDOoA7VBNQ5BLEr3Ysu3pQ9m+VSWaztSpdaJZHHkE
KmrXL4pIud8vUE+HrNu9D4QPRsCV9eJ6oM/B0mb5unbnXbyBkmbnER6s3W+HSfVu
Tf0wo61WkB4uAUjgKhP+lGOJVCoaPxhl5uFbRvueiAMbj3+Ze6dLz2E59s1GVaBa
aqUKCQ0dNuvKepkteDxzqLpJalwACjONzK/YbZYM1u6Bo89gDLB97m+i8mBSaFdo
vG1sZpzDGqqt5Y9lA7qqRzHWIhAWyLMBU6swqMUjbcLkRrebxRD5cv+LM+cc/veM
NbYEtxXe9p2LlGtw5up/rFieA5zRoAn1LhLz/tdgaTFbCSas7hGc1u+hiHv6wwLF
7uxwRtlh514ioYAuCGr9ewhzSCgSJQPj2USUP2iASXcV4lrKbDTPjefXPffauFTE
CI3LtLhvfY41Fmlt/sBd1+IV4lW/ljOc2pD9Im5zJZfk5/n305/sQpzUw8aS5VFr
7y4XjfxDXpVtSJNmcg7uEBll2D3JhU7ujiSyJaxlr74Cv+F21wBTOunO4lf/k0nl
Sqlz5g+jl5SVcg4qQ38Jq0gP36o3jKZkcm6T8+a7yr6LrLaRMxb5+OfKx5Ft8mnq
ozq88feoVJBWVjYC6AJk2ZPLcG6ejzlsVL6qght0PA6Qbs+pN/4memrBOtdysu6l
uFKQUg9h2yqjmPlsx2b0bIBzBiz802uL3tizJa+jr4qsFFWVDYD27FEoT5uwdwsZ
OgihqXtRp6n5gwcVBfhw/x6Pq5j0LXINf9DaMvsz49jVhhNG3tVNSYBIn0mSl93Q
YWhxNZRr17HAxy7ZglsBNWUD1ikPPHKwqDiM0HJ2M1ThFq1CKH5UxSPQz5w6XWhA
tLe9LuWvjSAij2AfYkZhFijpNjLqt8khbj2s0O82Cb/jHjzNt2KHe73z3oTfGxpe
48edZ+LiXaejSfvJqEl+Lm2ga+/N0w4Z0csx2Xbw1bZa7MwHONqyk4ks6lPT6Uzn
+k4+NGMfME4dPDMCGGywb5/iH+g48XOBb89Z6/ayzruU9WedlIua1Zmy397Sd7PB
WEUhI0eHG6K/22hLob9M/x354fM7yZLVMDxSyNKgLJ/2VQrrKUpv15eQhtgQiapS
nKx+ecDWGpsWuCoYrzYbJkSqH+hHsaQ9PNBurHLe3WJM6VpA9hl12wu4r/ude421
nljUIHQb/7/5ARXVb4SaKtEs6TuPoV075l3lV+O+fYjtjIId88GE1KnKmdFvuycp
M0dMSsKyCPR+8fdssqTKyTamzyEv/SI+0VB19CWh3GXLvFrz+GdCY5MqaCAHABK8
1qjG86F4SnHj3XqoK7aXvhNhGWVvZgKj3a2P+Oy7WSvGK80sET6DkDnDIdv2XzrL
t00NEU6XWLgZM3TB7bEZHmfEUiSsjQNjiDpxF3HsMLZEg39GidrswTbC8qy1EZ18
Xge8UAoLaZxEnPoavdaqm7Ap2MvHYttWNijvTxMszHrczfPDfOFuYRvVySnVQUMZ
fkJbC17KP9pztU2IE0uwhvDkJQuxqC3uZZzVLg0wJxqUnFf7BQVTbmi9iNIzTnDV
kZyAhToIzlwjWYwK5mqsHj4F5gni0HQevXULFx06F1zuL5UQvMh55UFgsIH7/7ik
bVJ3bhIpIjYVOHgqiiM/IcsLDuezpcFWvx2d5ZQJfIme7MdZhk1661uf7nlOif7z
nA7pUtL/P8ZLlsz+dq53bTvckErMMhsR+tmMna1U3/+Mx6QNW09FtptDVMrdHbyb
2vQCX/JrbaznsrsRav8k399Xh5a9kog9hizYqBIXGSMW1bqu3dyk67TNSie2kYHG
9zh4VEtcOHUr1292cEQc//vnuZiJnpcv6VpB748x3bm0yVvBbib6g9TQ3Y+s9xl8
nUq/LfhcXkY5JwyMT8zbsBU7BuE8/f59sCAweDy5ENuER26Tn5rJpBx6nC2kKCYY
d8QI7oQUyCEsv07fgvjQTNZdxG5qNB5ibTu3cJmTlcBpDJeaFhjPLh6ciPBS2lM3
3jb/t0HipPamw/CShWGi7+xFqW2jJpZBaNifGv/d+vH2yjsK5vRA7pU5xyMJ7loJ
d1YoXMG14o+uuJLUxr1nPMei0dnU4xDm7lJWXW3HXO47WmV1wBxPiY+jMsrZuj65
QsnwJCA/v77jEFTSTXNbgr2E3LgX/zunusIgCWAiHAXO0SEUgBHn0gSEqnLAMTFx
Sxevpsrm5YhFQTQ6dG6KbJf54IMs1IhOJEtdSXyQzyQnGMBkgH1bGl+RvbbBbZNR
5nqZdcYb2GSVk+/weBVwZGjjh6bJQ+eY42yf4L5WV5+KkXIjrz8WySvkmS4/aMXN
94D8cTL5y9nKR2VaeyM9SPCkVj4Q0cdDm/D8qeKyOQcw2QqSwNJuyxuqR0BkfQMZ
SW3oC2t7BHoqXg7J5d8FTnzZgiRbx6jmsy8Fj4Wlwl1q9DpIQgTQt9j3DJDVVHYF
CXKDywf5hQQzTs5Wwye/CsYjHKl9V4HkTf2Wy6Zia9oGHxpYPFlSlrToO4i8LPRe
vzfWqA0XWUfbweVoPyIq4rnGFapDmVr8Sk1XdTn4xzt7TD+SQ32Etbs3oIBpYNqP
ltkOFf72tpe7U3sxhc4Q3cmoGzcL7T3+yW5qeEWgOhNIu/b8y4jMwXgwAXNwyy5H
G6CNkAKVpFlYDRmJuvACFxoT+/yZ7X8kSffNcLKFIY/1/ankI6GXVY4InBaGQRQd
S15CIFblCfZXFk7LhAoX0SDTuBJi0ExLfd5lxu7nm3X1goBMA0NPAayJfWdaJUds
9B5fVEPfLIzyW7NDDaK71Q7U5reBqJWGKWqf/BqhcU8Bwvl+A/V22O77HSzgLjKD
fyImTOJD/g0JcOiBtpme4PpmP8IN5RiI9KNx/FeK/EE0zzsx6Tu23bZURcLWg6ZM
oI1jX+ccoIIfVjx43fqbm7Dt0+YZq0vkLr0RYdMrRuFZC6pYGo31VqK6yXoeyvrJ
bzF0JkoKmyOUNF6S/IEKzX26+j28C4egk+NU1LlzJ6ivHfKjxvHLfBE4i5T43aZi
2JOgEn59RnUZy0jFQbnvR0DwCEaXfssu7fc/KCWPGPSxe3dIGlcV0nufyD9Gt42Y
Sz0FV/7rw29CyZYjfnxdZr0fNO+4kK46/6Pk2n0/Ohoy9bnoTUgL92d3UHPmDFKk
1mtPZ/XDTT0+h2K8dN9uwcxMxeyppGX/UNu8ajPSY/lfLpvzmpk64pC4GSWCw+86
DW1Ty52zIoo2ZkvkeEHSRV0SXXKTcpW54v66GXXurg/cL/H55+tF9Urgt2U+dDe8
vOBKdjwkWtVvncbjQL4lAENhRtMcy2IlayomDfaBGwvQoR5wMIlg/Ew95QPWnaGW
mx+pMo/JbNlWRcsJpwcWMrgRV0fclw2N1u+0nPyKSjJH7unSW20oc6lckYoy8Gv5
9oPn+D7QWPXAAdCLMzoA6aJU2GXOdvWsODVFn+M5AHVLDmD6F9s4bupXZXZu4mtz
diTeuBeoT14gS+/cBxcYgs9BtYDGNGmbiIdv3J0tSs+9j9NMl3VpofQV5LA4THNY
0vhQ7cPrISm6xGyAf/YHlTqwEA3nOZb+HsfyZLi6wyrw6l0FHZ0BzV6kdiY/G+2V
E8BMfZOQ549irVGg8t+CRrcgDYRAZtt44y57kpIr//FYkl3QjdiKtQ3Ganh8KNng
rcWRuhSI7nfdnz4DbAllRCLQ6dcwKdvl3tS2vbnKFP5FlfU73MPPr0jVMHk1JiRu
8DwKviSIdAFuXjSBR+06BYDBuVHNmV0eHB25sydukwWrwto4DKLt15cUrfnATImH
lC/FBxI4uyrlGv6qsSRrwJR7LMc0wL2fAiQ2EzMteGIavnid/aZT0nwzn5Tj1Ixq
JCjj57rmczD3q3EpRSug4xvkvYmNGE4H1ft5ENylFbdmCA/+2IdhnccMRtW4jLeO
eIeMA3X0oMY3Jiy5U8ElXbs8yWuEj/HHqF3hB0DntD9AVVthh1WYXa/mBeFtBX9y
4H/VrKGWRq/hvWrDRYn7S+b/obUjiladqRzu2BMDaX/upPGLbvZnXkH4lo8WuqnD
W08YNtsAg15yA+7v+XOAWp3GfdmAp6jF7FdQ5NIzwh+wVopJ1OILpZkGYhj8ngVk
YgvY4dgbzXhSFn5U8mTHPo6IeQIS/Bc07tAv8Tw0FIBE0JT5mmHnV7sQrEjKRk0o
w/kTllBoVOYfmL7voICQ8n/nuHxjxg6ZI30KDnjzHZ+gBFCeW52ND0NbfX/o+85n
CuB9bO356PXFa3GhuqlblMPEXJDEaJQlyh9kGTH07AdJxGVaVyXQsWuvbw7V3fB5
uMHjknnCyjpnVHKoIxZDqRUN4sBVfiC5xNNcre4ZS628Nuc9VfuSC48Su2PZFyd5
UWPPfVvLv369iYlKQcxZK3Lj7VZvI8qllPmi6hwA+j+mVdJYm+o6TtRq3VFHNySE
fXphERj6rKnmOaOTpB9rPIjZilvRvA6xcE2qYlkTNB0t1kGv8HwKPFLKTxW3WaWQ
PRbfDz1Ljj2UR0+VdW0QDgcCsE74E12IDkEtMXw129KwxjU0/PPFfBTjDBG0lMaT
kDYQvsLsLpqhW99GQMhnWcnemb69JvqIgmOpI4nmcS4Mb3JGlxFVwIGMq5noeNox
gNRAkRPK3HxPkMmpGSzWo+Do2U3+kbKsKfnsTQZKWdSjqHJ1Lfp9euB4MVC4Fzik
HCTR73Tnz3LbazcACCyzVXy/+8OR5TblxUjKJVFWSjFTcGXnTzYzDGRhYH/YdBUD
7uNiq2/5nAogEj99qbFi10EsbOEe3knr0CqsuKtXMhF+4zsYAmaObIOzlvMytkgc
FD+mfwrWz9jNXQTtOiYlD4E5ozDW7PX6wnlD0jqt/m7gi/75AihwMvh2Zu+EGV5I
Zh0FU/jTaKGozN23Q46dWT337VRx0uZBlWVd/fTsTw/d59SlFFFjTlkiRuuGIgND
R3wj7dzRKsMb4rYvGoc5stPrELJTtyATNrXPGWC1EKPTIZfkRwAXlysNWf57KyUi
4c3HyREvCWh8GM7PRrltQfJRgh5Ik+x5aW26+5wetMM8UCQ+lN2MnP07bzOlyGyG
wwttOV05trDc+2AeVl2oLO9OBS6lZFFZ3VDLy2J5w0bVsVBf22PfsqnfijlUrRLM
oQ2twAhqKN8bBydXZVM9UML+5cNTQkAuUt07sb/TwCTy9xPwiYJo23OEO7KpdQkF
/j8KZD2BLZUOcCQi6pHzn+cvsDjqUFwTFoXr4KuRfSzeJ8J3MCV3qJ5LQi0hXZuF
ls3Y2Q2pZRrHrIDPSuJzMvl6IT5R4GKTz/OtLVqnqc4CB+paDCnFtjk9tDF5vvfI
Ao5QpTAzrIfTnrm/zJtkoS/ZqULIr4buvovDWN7ecFUiKU/63BtnY8A8Cv4tH4lg
d3mOOf6/q3Pk62lIhV9dlmkWkvRGDx221UyXzbZCdKx/t+ZUalLInGGrhOKCtuSM
zqhc8x/hNo5b+1jLF6BphzrSAfnWGoo7Z2lhavTv1Vs4xnV0yU6REHhhgJd3u6K+
D9Ma9xYeIE/x1cFJlA0NoAo19rfeKWg3yemrFf7CIYhQLDTXygndfou2cjRVJxMr
XcwdXegxxuxqImRCjgzS1PrgFFiHgFwwnESA1A8ZN7ssXxf7nFDBpwXcwRwuRv5K
paaBSHH0Sc7tzPAfiZtfyGqeYkvA/4JGygibMQ6HloZfVRFupljGSNb2ZEmPYPB5
ki0is/QKJhRD5GWVUZQriWM3UNF4jte4knQvXQTw0PRw2ptMJuvPisvlxoXQdjRp
f5wT/40YNbuFo9zrvVZ/kv8SunZS4BJw3p5VCu8cgrgsY8laze5YE7V+1d/38TD+
EAsXOiiviTSJbUxNKl2ekAEnvVL5o7iykIc7bCuLkpigA1cnDD5rCRtDYE4RSPiY
U1kjme+RLE6OtF6q7xK3L6BEroyxybLBkvcPXFflmi79XKJqt5OAGDZwRdaNOCBY
fpvPZ8fTVUmQOI5tcY4B7f/hL07yZTmvGC1YqJhcBQrDf4w/3NzFu6WEpHpUKf8g
b/c68ZRy/kU8oamTc/dx/4ZCW7vWCSjlBSarFb+Z4452pNvb/ITRQV8unZFEhtYW
tn3I2looLoiJpBij4MWFptlliHt8Lb02piRM5DFtHnxihVB33Y6aL9m6LAs6aQb2
OFBRzRIbXBB1WszxvgGTsTnpzzrKHPJ15NnYUEtxT0RGPg0tKByBYGMaQqtRlKP6
mGkIr0FK00Wil+jkY2MVLoUJs456MPIgxrxaKLPNTM9UAnrwp+6aaDwpl1TfmiMM
DkMToUxxYpMEcligUPJeFVCTdGJNLWFLaFW+gfqRK39ViIBlhWRXsSo3ejfOZIVp
9YzvTldHOJipcsLI3pdAPhjRDtp1Jdk1M/u7d09LyxzwX38y5z+Tx2Xd1USAPDCl
niZNIxYBLVank+u4KymgFtyxB+xUel/IUjvLw2wpaVR02pwIX5oWPCOjUgKtogQm
6zqbmUfBElx1B+9TaC+OUAlFZSaaurqk4AwKgevOFGSWrIgy6WQGPJV5EZ2OrGfe
Ix9tgQdUn84vFzpFLtQlxZ1qJMix5HiOJ+ATSzgFvjJnnKywfQ6n9DP3sCWBvVYB
tlTAVAui3sjzPJJSd52iiGb9Saf1cnE86t3j4/wjyDKgLQp8gwsQ3FrOtSyGvpsl
ts/+MehHmGaj8nOQOu3Smg4G2e97EPH3TRLZJxXS/oJfZE0EZbAANZTElQE0pRN8
bU81fRFkl4817kEpXHqXw0ZpiQhaRommbDTxlmN4mq9CDHuWbmxIAEC/3pFuoEKy
f/+jJ0klzhbj7YsA3mhwMPrIkS3xXWv368GaJh4hRAUufzQj2/m3FL7i8Deu7NEz
wggqAFsfLh8YEU8YnoO1orE+rqTFsN+WqlNeoWGDcbiLKmO1Q2gbtiCebzNF76qK
hQCQMkM9Ck/Ce+Rqu/6cTA3UY3dsHZHfQD+nb0tTM61fdsBOmNIyTmTCfpF/ptgm
7lefNCjdgQ/uQuZSPdJaHVDz2DKz0BZPt1BpWOsRn4xk19ncKxrEXn6LdtgJ81oV
YNf5tB73cXe1s84zh5VTT3IpNrNmWli8AUxQZA7LoZT27gVuUa/A599MpCMRb7Qd
f/mqIn+tMbzp4ySZAjXB8url4MYR0d5VuUnJm+8eyF/FwvzqXgwmqO0/X800kPmP
cBS5DgexKI1BM/RHz/E+VZrHvDp9cPPnEwyRqZf8kZb7IJLU0FMw6OMbeAcVLr4y
um1hHFWZve08TOnTWyFVZjqte7Tq/y+jewdZs7DnyzMkD/QNbbaXv2SJ1CgvtAdi
6I+lkRyqjppyb/+FnJ40OSvfQBynnTPXQszQj1aYxxcFA1QKuqW8X3NTFkJYyywd
Nz4wuEi8BjAJ/9FAVY2L6+re6mNo6yAveNTzw7o06Kog8GLAyIjV3/lVNBolrDo7
+phFj96W0qmpYh4ocYtC644DIUyLIPqs+Nvf1QkoRnKvxH27wBCCiusFiby6ALxu
8FRx2tzolWE1WE+z0cHLlKfBCWxwfr9J+9ORBYEjH9o7T3UphEtFKt3n0dmGJ4+P
JjJzlTqw8VOvXbv6eYS29/0GIcFq7nErlOc118hWU3tahukwUJUbR/fRkFA/hons
DwrIw/Iujj6kbrtypFrS/F7iZK+5Z/0AdJnb0nAcMW09+KUErTfDCbz89KlGfhkV
tp+q3SMxOV/nF0PFlQta0t6C0HDDKTp6cwL4phiWPEBBw2BK2vdp4Q3GBlvWFH2q
ZN5FE+E7A0pHmQd62CrehS1gkhUCipx1OdvL1i2zvzihXOdtPCvtF2H3BsPuKI3D
Y468LTceA+S1aD7yOSdXA5rq2TaGdqB1i9Sl2kYSqRy+YgrFJPABNU6apCxba2O8
n/9q7hQk2qV9MxINszbBEqJL+PZcV/ZTdXhyzKfwzkoiMFbt+EC3y2XO3+cOs/Z/
qmEAo9enKKrRUsw8Ej4EZ/AGBwEREHPyRBEBU+k0V4g/37mlZYM06+7bsJpZbeKT
+as9az3X4AugBfyYPkqXgVbOyB900hBwUp0fZsPXfPBIrxVq6c+cNtm6iB4Ck6N0
+uBRbsxAsnVDFlLfmAIttAZZAbUS4Vxf5lPYozT+fKMmgenmjDb0P9xQTLLSCIgt
t9JfW0XG1N9/0t2A1NWntsUgObk96ajGGZ8yA9OXD/tU0ATXNxbgcWqUS+fYs757
9NVPnvmmUfqBJh2YeWxC5UHRv597g0Ux8zOGDOK9dOIxJNNeA9rRBoPjGEKaZSY8
1QVAlZUIc6Tkb811Csf4ft28jPmopu5MPWeiKPo7qqV0d7IKODM776W+Hao0WTzc
utDQqWbnARYVtDPeMMnLf5eKIaSY97TQzclmDRszTo52+3Zt3kNG5iaTsjs4IW5P
1KYWvenJq9ObdLP3iFP57mWX/uLLNDZKAoAFTjR7TyVwrYCmixsBACu9iIPGMRmf
QqWbK2hz7D8mx9UkfECiYum7V1DilyO6j+UrrIB0l5TN4EsJkf/Gy8RCAYP3eOLu
YFQEy7sSwzv5um2Kv35gXyPr2c1dhNCLKCUprVsdvK6m0bTwtDQsxfZvGtRgeJde
cNj5nKt33WQ5tg+BKHcrAH1YdMl1cIkSx31mu63DtIl/qxzZ8H/hzkZoOXNKqlcg
WdnYxNlYrxgqPAKPnRVSqHNbNvSnnLMQ0RQuj9e/DZxlrhJ9dUV98gJEQJzF7+Yz
aXBV4NTzqqmff1sQMv2+W688YThXZU8nW0XHy8eOGQYamb1iA55KDkynEobddEAl
fzPnZeTH83vJqZwwunj6JnAqsIUP7TILNkpkv7ht5yrnGO6sLF5/BB2zDTNMX+bx
ehEPjWDdT/movtddmFKU0uTxS7XC2JE5ph6cEOAc8Gs5fkV3SSga36KE8oBsd3zv
0piyybOi3zcHmZm1MudLEWbisUbRDC0ih/RiPUo1yyW/PV5bUk478x4p8hMtWzmS
v8Z8pX5aKxSBhcDERGgrT0iQN8dedCTJM+ngvx6kBtIl4iDXYRN//V41lWVe6lQe
LrtNS+Nx8+Ug2LMyFamZKMWou1htoQo+upsktOspctnGKcWSBwM6wr6r96ZCf+13
l/VQ1GGBNuNlhyE+p1Tqgck5u8joqv7/ROrLaToI1LSaYd+P8iHlS3CNmpY83r4A
l1zmwDWsb08mcsLfU+d9PCHmsBFIP1bZkmDIFfflZE5jNVcL5fkq9EgGERmL/Ds3
owZDn1bA29qjSsfbToIdJX6XspTl7dEtU2JQguh6MSschi3oLL2sxiSk2IKCh+fp
UZoVck1rA0oO1uKSYdJXJ7dWuJsi4Ji0+iRvJ9EVgKT448qA6kNkSfmq6yMHuqKQ
UxYGDiVJKOMGb0jaXSc/sN7x+l+t70p7M0dfszXGon9yyp37AmeQtzH7M9Rn3Ij2
UoW+w8G8YdBGPTSZs1ckKaREWw+FjKFkQgJSjej+6kMlG8C/qfSd+m1zjVT/leDF
DNGRPQEcA5rR3UbVEeLYNux4x33lynYtFAeCDyyM8lTBwfw7mM75MZB4j1Q+8Ujd
fbD/vCwQmgA4KBl5EcZiXM0Tse0HtNHuIilrKPjGV4OQg1mqyYcT67quj2KvL5op
D1j9Pfb8ZfKIIFL65apFnnLsAsi+Jg1wmnOZdmc1VIWnQ19Wt4u6KRuCeDIeidKw
TW4tQ22RRB8bNMjMyZJv83I3dmaqLSGDmaUWWn1fkH10LX/x+sXCv8NW+AXx2lGn
JY9eLnDIZ1llPJOxyQ0a9SGUHCRDvoIDZr83vhQJN4YbdmC6it9WwEPhnrk5Vacu
o8OpWT3m2hxqxS181BCStIoAYEQnbt1Q9bwsBdIbEpXc45oCSl94RVOhZYwQ4E1+
m3YtTV+ornQJ7A1FSliMGqC/2gHR1mkoCw/4gWZ0Y5WTcVwMqBt0X8+GmDoykWEa
MGSXaIy5bYBMFU0ixylGRo5tSd9TnR/BR0zBwn0QKa/hglogfOTMA2lrdAHLo+pk
nabZT4ZYldiU6UMThP24sHjeuJThQ87jwA/zoNCNTJu4cTRSKhhCMpjTzYuIdN67
pl4urnVnKV2GzDNwoQ1jPYn7K0Uj3kB9JUEvz4kfKiKnnj9cCINQKVeJ8kprZWcM
xRNnxiYh5oCxJzXIBdSm1qDuyukp+FO1gY8gdTqhv3xSVCq0aSXOKe1XpCk/aHC1
r6ouHpNgg95khyufwH8ANhWJc+r6DO78ESkrl4/iNbc2WSAXgG3q4jC+sq+CMIEg
fajhWmUFqY2je8oevEqSi9jBh66fqo6UmmjLRUnzIIsH84AycrMKMW2kpBdZhU46
M+LSiFLi9jEbvFMc8TrgIEs7Y3rg//xZyGcqx0AkqfvLU5SlGdIK+XREdLdachNt
Es/GUtlWlFv3aifg3kc4MByPFoS+jTNPVSt9pCtopF5bL2YxLvyre6v2vXkzEI5D
/YuM30FYJwfoHqP4dK2qRpEs7FkdsIG32t3aDHSXaSpa99WkCHq7U/xwhESfcfmN
WQQT2ZaiRQEDgAmMcBatN1QEKZK9njjuUz1uzD8z7n1PPid76TmG5bu7OYjdRZgv
OPrkMHUqGFW1oVIdsE/IFy1ovScf3iFHHV9Sa+QE7Ll/joPTVDuXvIxvx3h9+nLR
yoOwUU1xonT0ZnaIMm1kAwj76SyarkU9f5pM7RC5Z5YM3TN7I7hQaIjwXQNYqGZ8
oVL2LLESp3K2b0LWTTOmEHH1UjRdJ5rK/AOGt3dtn3ODCgnWXbwpbJ40KhYLdRGi
0CKZ9WQNpVCvGso7gh/wYd+rJN8XxqpHX8o9rMKvX+UaaG3C2OuYOCerTPHmiVxd
TIoEPCC6TuIneuFwiqAzshuHp91JWWuGW5HJyCRr+wqzuhdN/FOLALqKO5wHm0Cp
R39SYYFZINdGmMNDrJpRT/mjrmR5lwB3BS1JpwCpSEwv4sDKqbb61CgqSVbCsj25
nbDFvnDFIOr8mflQIRih8MSja5Uj+ILaIWN2awgGPeSOOsLqHIttzESydNJIb85S
NDPm8QrHCN1kVAhjz23fcpnTT8kENNZEu55XpNOvWX6EogQiaecaYVG4n33VgW+z
AzZ/P4KP1VNXw0jfU4++ixDHYEGXLu6/0Ld1vMMWOgZCMJV6K6x2H3a2laMNoSb1
nB9+HiWnoJAS2/eGG71lK0Bps1NGncxjwLhtGxIPA7QD79syHnmFHJhVXwm1SFU0
RtmXSHmkxR4F/peGlKATEfnj5wXbY0yECZf+7lQpQWsiz31T62IXJqQWiZP49Bjb
6TmLsed+l2VbaiuNrQ5mhc3V7wxphBLNWiPLnosNkHNDZVTXt5Y7QEwEgGPZBQhp
lIrlEUcqp/uerLkcZnxR8+qOqCBphI7DiR3nY9dHAe5kWm694bUZ+7GgARu/Ch0V
boqutVIOBBzqYA7wcZt7/cE+TGeO7G2hFbHWY5Kv1ipOg//vngPv23ORJ/crOTcQ
aptJgygMamktjqpv550e7JnQoB2+IsFD3PI466oQTyPY4ulv6CJIEHgw4ixFhEvf
L8DdGly6jGmrIs86PtwbB4wv/slgy6xQa9uoczocp6ptC4n2TqLIOygpBCuHn6J6
NV50lvLLbw65BkUcalpX+f+C03Xn4ODBD4/fMlRtnNyg9TLg4aYtJD7QaMCuS0p2
yPRNj7G5f97BXNUNTqYemvxm2rssmWxvogOvTs8l3kbteqEwpD00Fi+fgsDzHR+s
N56dFWpAL/yk5hcku4AAunknAwm79fCpTACf3fdWy3ycrSw0NktBQrI7GLYrRVin
CStBv03jrOdBiA0lKavTax0MYyw/8cbCuVPT8L7bRTu3KSIvstx2W9F509BrlVFt
h70sYJULj4CDc/ze7xDnpTrfhkNRecIU+v7rYdzpUDDphrEsHEdZ9MbW3EcdwA2y
5pS5JJFS+EJ/oi9usRJbjV5HbpEnBux0Rz3AE4+ksUfX1umhxCKzAst52tEDGF68
wz+OB64jT0RPB5xpMjj6W8969FvMgrW+XfVSuCL60VUfmXcp50+2dPRATwBrM7f5
jCJlryLzxZfbSTMRD/jCbRn3UW5Lsgc2tOQn/sZ4FyB/JBaVh8MIOC9vKp5ds3sG
evdtYwQTs2yck2mtzNcAt9ZEOndvw3yjBM8srEzvwwcRpKcCC2qMkcGfGlhdhTVd
x+u39OVXyHPElBM6OxC9PLUjifjMqJtse/j9Brwa/HaDrvpDAtVpXqtt5i7xm0tT
uINy4UJ+SjDOXLqs//dQwRtPYsqLNKdGze9zbBuSVPVdb9c7LRNkFutTukEpoIIg
o2RYWURMVUM/JG2CuPtHK1iMwuecqF2qdLkheEVBDXYW85tfWM5EmgsB/NLRIAX4
IB9wPUxvatewSZwA9oIr7+Y+aYx97zNXs6pFf/MJ3DwS4dHVfXh5BD3yXhrlK8AV
qjCnKYW/w9Xa9i0B2CPLWAjuEdI0X45oIWn3hpbkzqSg/n7nI6j1cGxWq3zvTHai
S/BShXvpmG9j40z0bcNK0F474QA8YAmwB+0qw++qH3goUDqo2eR0LOqEXE4gxgpJ
gWmvnTCnPNVTVE+RA5kJm74ruJPPkXrB9kK+F026AOLfVXrwovPdXuJggYdDnX2u
WdfVVs4D9if/B2luWsWKZ2HZwn08lYx6gCg/QL3nBi3GBLVZ0B6RgXzakoC/thZ7
PZ3NtLwr3yk+UHJCwDo5o/0ZCaCgYjsinNfxWAnOTE+Y7eSsL34Smeu6t4SS/+aa
8ccwxhk4Eoe8xZggUDWi8WetDvIjwzB7N/N3s7NynGWVQZNFJ7E4FmXgd+ll44jH
xjS4vvsl5lOaj4UeDkvzUPoVVW5vAjJaXhN2sAKeeQgcVukJ445jFDfah6+moi0I
oxzuj6JOZPPveK5adZF9+A5XKujZB2q/2uns4EBEzT9SN8hDF47+k8hMN+HJn4hp
L5u6pS2YcgD/Gbx87A6ccI3VTvlylk0qMes3bhB+C1JT+Kgcvk++us25570RY4ag
nBnZqEckGy6Kh3/UMQ08TPKdNpmHrLwo6i3kmFzyP7FMcQQ3+tS6BqD3Bhja83M2
u38FPDx37R1uVEMK5UCY1hVoWl1ZgvF2f/dlg/2ukW2Zdt3PRl2+fM0x7uCgnN+x
6iM8h4A56+JU2rccZk83OFOP6ymzXTgWKHaWM19AUCincU61LV1t8NwD9Fbci3vg
UQZV9SR8JMApN8q4ussQwd7g0HDLHBssLfZSNbypvPw6TjLxMHkR3UhEUnlD8GV2
0SM6b5Q0XJ/TALEleUVYtutzKPKXT8O+2U3cEizX7pj9mgSBVVNWX3+F/PiG9cg7
LmBxw2hj//VohmKljSi7c38Rf2DuxYeGuf0xfeBZSwTCpBJEA70Y3u+EsOPglozq
ztcN54BqM4ogUKWPt1T6LIfbSPC0B1iBXSOV+WulpSDM5oSXL9fiLqLznp9UYbjz
FktG1sbW5CeDn2cuNLzxfhSff05JT0HRDizBt53GhY+BWE8C4GXIYD5fLrga/FEN
7yZ9XN99hyIvfhbhFdpITCzqOpBrjFPHDw9le8FJ+5f2hObAMOejr5W/n045Y5XC
YTQJ5nVeRYQXUi6ntAm+uBmNmB3GGuJ3nPXOy/+UmZ+jEsMMLC/t0onDzDuPPHiJ
CawdrakARyl61Z3iIA7+/bGaK1IcvKp4qZBzBxSWnLhALcphAGH/R0mcuyDshmDA
avD2dHgdd57zVEJkncQICCGznHTvDU4prt+fx6xJI3PxQulnzPLJilpftO54mGX+
YMlqPxPcUN1jF4TV7KeTjA8pFFEyFnhjHeD7gvZ0hzR5RwwhYutbtJ9iV7BcV6KE
jNlmRq+WL1ABW0Ay0uooeue++b0xzsy7tOjA78xByI22gEjuKFBoFEI4/G9ybYC/
hBscwizmC8ZwSRYBnm7THXZ9Vq79DlxL1KzaXogC7Rp2bymJEnBvj5j2vc/b3RvG
Mkj2j6dXVp5t57uUPka4AYmKf+ipOVT1nEFTMA9oM/+ULEUUFBiai3pmAmLAydl4
fIw8Tl515hcLUI8KtupMW51Wdr0ohOKbnVH9+7FgrbAn54QASQmaZtlukYoIbqHG
G+zc0ds8Bng8nbQQElI879herpJ1ZlMvHfY7D761AOzlMmXk8vsATndqNF5+bxnQ
vhHtFH/GWi4bsQCZjxszWqxpvl9RxEc+MPYrpxSlrEBAeDAz/pCTbc3I+QDpNdPE
9L4ndDGlvmYpDy4DMUfpQ/YXJTAGPMz0McgEeFGAj1mPb7hjwukZAMKAeWrlH5cJ
P35Aa29UTJXiQHQHhFP3y+PjFuh/1/rgXLVWRtALX2199bpwzWHZnBnj4YzyypBB
r9ZngasmJYdp9B44LL8GhsVDdqo4pJ0s+nax9THCTUP31OQjjDMk2A5PSWeYz4vP
ukWWsyeOvouCa35EU1t1PxZmi/cKQ7d9saLqJ56BpLz5z5R8wNXditNcqYbP59kZ
ECldnFxIKEEb20rKzXtPmQdMO3dqvZefkXjSi/znDBhTy0JMDwnnmOZE9fbQ+9Gq
fJpM5PCdOOwyzelAEds3HahQOpaitTWoVPs7OW0g+UC9G49NLpcoGnyHevojRcmP
NHMmHgzbXXEPWiPOhCDag/ujCsa8zsaTDSNA7w5Q7dlmOkj7ZxXm73yjNmD2ni+J
p5cgIZvf+5LcNGNHvlmzS3BxzQKI/AAJDz9IJBKJIvzfGzM487/xLdG2d7fpy/5T
zgU+OrMRz1UhPk2bcwermXTO6cUMP7OPUpWxHNopr1W3bL6f/12IZitqtiVup0Dd
Fw7VM+5ywaL9GOWI7nI3pj9zPAZL8pcfvZ0tokQ3hUFLRmmuq8wlowMk/u0dwAPQ
dqMx729dRWMwRBaI2paoZj1SorLzFK6GiNBqNmGQ6kO3LpnApwWydrqsrUI0HrTd
06mOEtNkOAlEmA69d5xHQP1gg57zNcwHPDCGji6fG3WIPnNd5Lt7RhMv+M0sBy8e
lXfVx4uTkrMwr3wLmwEac8+AgTpTPFlOb9Dtedff/IzOpN8QYGZtKehRut43YdGq
HIK/ORL2yDZYpjG5RU/7tX11QQiTJEk7g/1jXGgdXlNwnr3PD/Q0Zqa0k1EsILPT
UG83S2FSJnvsEu6WhZCXI33JF3eLmgmjoshroizukj9ctlFDNzeklBFDV4gfHUzV
HA5lK1Eggls4MSB1iK+/FdYlP4A97Ke+CPeNO9GAq95n6jxCqu6oFmAnIaU50PMJ
6O8PbHujchH8j+opkSNXXGlejg4t2bgvysM1wDYDmVL8IPn7138jGyvl2Qsumghz
h/Ad2dgZVG+0XiLP88MDARDx8RoCDqlzKVDeme6OVvQdZKwGDuzZc1XjctPQ+1fh
tAbyLIICBeMmYvgYXTDk28GS7yM3RvsTLnTmuMenP9TsQG+sRETfyr64UBoXB7fV
cCyFSH93QEPzkWT7kQ8D7SBCU9dycp6q/dJ/Xdlu2ofk3JiZLC/2kymmLxYCOi1D
ln9HGI+dXgrlLosFDXEZEMQ8mnPKx0s9EhGxSNjbgic7pJ64gQmv45K0Whszc8zt
/khmvhct4d6ESuSbyaHa+X8WLKPgSwqQTddvZakVvR1+xk04b2gmDnFR5O9JgDR0
p+nOkJDRr3FwjR9ADog9ZIAXkK1eHdXTqb6BzAQdBK7+w4lG1rrrBrQgTNhBNwcM
dXrON3eQHgxoY2Y887baNxCJ6qM7C2i6/JL84Zpew9lAjvtjVgRjxWgT1iQ6JH/0
qPuCv94Kjerw2TwdJa+UaxwjmQMEqKHaHYqxZotXMEoi3MvOfiGCShBiDM2+FG19
BNY+9oRcvtKAulXp64lX4GYnfTPe7raTf3bM7jroQl5yvDlNKXYYPMpso7NX8lk9
dNFtPelRdMdk2RFQgW0m+jyznFZ0AVJ7zW1LD07KrJT0KqvmoTBIS5usl+MvaQhx
9wtFcMi2VTnYFHM+SLbH1iWskTUZV8bU9H95cNPnwDzG56qKJbrSpLUbRersNRaR
f3qVf79aNNEUN6S6MDC5XNxA949lAFzm6m12hnS3WaxtTwGFlxIYlMuPOhG8T+TM
kousHwZC1qymQHkEwU8f1cE1S25et2AOcz18gMJrGxSITyGvTTK2yNeSdXsEJ+Pq
7zDg4d/AV6VRUWzo49vaAZGKtgrdrCDn4Dh7hPrJ1W0AENm5QvJdgy6761W8OnDV
9TCmdrxuyujNNAoB9cNBvGJx2SRNN3fcrc/DT9qRuifTPohv8TeCb9fLokGYU7BQ
prR3TOi4IRx5FincuMH736/5wuca5pRlgw/wsT24TktON/006XgXk4oKjO+lkOiT
+6j/yvWcM4N8KpGmWiVK71mrwb9ZoD2ONZ3sH884NDOfk+yTglT1zwx/YnMC63gS
3zVfaQ9KkWKnVROBlN7mXYz5YPhGE3MjJSR00mn5oC1o8NvT+2Vi9Pd0apN1hfZS
y9mu3F+WQUxBW6r1Q2aBtDiuRm9FvhzJYbjsPvIian7CMvsi6UkmDY/WXCl+VbYC
8tugtL57OE0Vumafhxdjo8uQ97AxjOQeKECK1V5TUfLhloxpC0t81pYAe/O5O7OQ
nUHPvJcrU+oBFLMR1j62StXSZ5gvgDuZAR/iSLne3D+ZwkvDqhVPCYxGk6XVJ4dr
RkDEF7XAmJFY4r9iGUBYMTGEOX4/AXCP0foHHveZmULG532Zi4CPJ8jvcSoCCNva
Agh0YR0HMF53y85fH+omC+EOD/iUkbyV8CzMssK6GKwrXU1kKUGQJuiXuU3HN+Ew
QRGLRhHoDASQTwEN8YXb7RA3Dq7QUJ6SYZLc9Udq8Rxcg0vI+p3wDNKK577N5QJL
Fz+4ltdkzNNpt5r3e9S0ddyzO+jjBJZ9Awbo3criQKY70zRqgJHHJIV1oJ50ofB2
BNGtC/Flfu6CXjfqcDKbT69f2y2WTF1wX/htc5vgzmWTxvqBdEmygy+QNShCWg+A
TqSjd2JoQHmi3ghVmn3syBD/1YckdIKR46yymxAN1GSMYo34lyFsIaAJ7cTeU5ct
iHSrxnc98jHrOYNcMgAirrpqNZDjHux64wnVaO6cB4cKHeaqPWyeNDpOU8qpAfN4
iA04yvcgbvzJmKdGO4g2fG5YkyIMI4ZjP3OWb/CM71lbHv/v8mi4o6inOq9r2tDr
PoAoCgde4lXEZmxxeL6gD2j6P3itxnPmOiz7Ztk4r4mYHQYBv50Q3hILjcFD+6Ip
A7lYf/9pUfrmJgLFsOqikPHUkwlVH+Vo8BpFhUISBIwWTbdnHp0MWmmXwPw9lCZJ
LtYkr+pFX5HvmUryCap/9LeYEYQdgpg/zNqXLX/GnV8TbBSzNGR9S2zYYmKRhyNq
rc3+MsTUNOvO8VTRxuNQ0aj8ylehs1sKeSaeUNiqMhd6P+emlwN9wxl9QC57oPB/
Av7I8HOF7Ho+5xv6oX+1mW6qTw79AiTP4FdlkPiT0Peq/bPpTBCNUJ30rsd/+vIE
OeWaYzmgczqdE71Lq8R7F4eNp0bGi5bJtI5dIVTkkE43Txt9m248ZlTMynaw4OAl
qwJnQegzMNh4DXe7rHIRCt/aGpPGBNQy9IaUvYh8qR+M4zTRhICrahq7jCQ9JfZ7
xWNqSr/ZZVXIdvTXodbWhp6dwmnodo4qej55tBrYAu6tOOZOhmcJK31shTdiqW7c
0EAavMbKGDINobRvto1HHNACgsk3YWSUPGIoMdTPCLt+Bn1CoVhVcvSDjiMLUWI+
a69Vw05mNH26wJYuI9ACEZeusm79HMM37+zBND3cWAj12kGRHMngRxqs0S1rwcNc
3fqfZeMggMO00KbG9nt6nxJrYxtMyww99w9ne0uvcA7iFW7UBwqDGa0rNcHt7uZA
rtK6Uzc5uyiRdMsvBRchRDXATOKo7POuJf8wkc44zCGpxZywWccSLDSeHuvfyKlI
orBRmNJj3zcLIZS4469pR/zMsitxUDjRMRSalPAxgMxTRsu7agU3SX0GZSsn0WVA
k4bssa3G+aXdn9MRP1zjxH4vUn6P+iibWA+MurNt2ebsOJ/mSB9MfF9zBwvEvwrp
Y1/icO/zLmnB0DhhLRy748C9o8mQRrHrwETG8l+byGjvWtBFE0C5KewHTYKDJiHY
NDNsGV5xllRSpmPaADhy316KpBY0Ii9zbFq0bQN+q3u8dosC/Zo7GBTCIUsbqzcr
gMYQ952p6fwr3yXDspsDm6hM2x1eGqwx8Z0QdGGgIcmF0dq6iFflO7jakL2FbIcp
k/mmGOsZbZqUrP0dfh2fJkkfVdklqGkJtvkDoMKtoME5639rXr9sSPIaW9dAfAqa
9nizpEIr3HDSjBCcpZYwHWY/2Kd6bxs1sfWRlKH/HJP1ySLFwFtpj7zUImsrBgjx
IYzkgjlm1R2P+ffJN2ejrHwyFN6khaQr5CI6FC9b9EUBDtz/yEn4QWqM5CniP03t
U7YHdFiz0PEDHuZ1IspQpIb5D6aB9jlfq9lsspG8xxVrzGX3G4GUtIjLH0DMzYBY
Y/akYZ3eCEnf6abjBKb/YkIuECPzPSn/AS0mhLFifLCHykwDhFMip+MB2ABVJjKQ
2VvVNErxq+58uoBYgfk9bxzalqXbhfb96/lYB3J2kuGIAlQuOntGFTx2kmKg+/Md
NRIZ1wM4jA873PopNzih1jQmzehuN3STY3nJZZmcju58cbTz1Y7NgajoVY4s+5St
O59U3eQB89o5h1zjiIbCwGlKhaiJSvoTJCSqEQWs0EZzkL9ry96wIElE/LNQzIUT
1Ageiiu2IAw5HRCmjVKTqtcQu5A+C5NxGxNjLoZdOJztTnvDJmuc+00dYgaSyilW
XGo4Hmi52UBj3AlvTZb4aGxRvxMdlUOqEEtP1otMezqtKZ33NrkszDnAbaXCGiCG
b9BjRMqN9+PjzQINUqSBiHmKKA7dO+nfYl0UoJWl05zLbqXZWJJJTZ21HuuU4CSJ
/YJjG/deoQy1uRssniRisX8XkZITkIX9ZzDMqv5kSWdEslWvENpDNV+Fp6unLCK7
Ul9/brTPcnLDW/2+3jXMR/GwdH7nBQ7C6hygUdWm8gog2ErPHuH1pwVcV8QiYMTY
Ix/9O0GllsizpDSc6b3APjRqtjHBqa49uWQAoQTBOKzdAB4LqLVt0glJo4dLyi6E
nVX2tBTeGK4nQYgC9mIE3lsqPu6SKFP2MnOLveflBxM1A+XisabLuYR0JTpwCboQ
FzSRalfY9TJBfKl3IITAtGsZphTreqtabxVgNSpGZ9LqpDVanOUsLEeXkmUokkWC
xy2d3tQSu6+B6keGeUh8HxTAqRM86MS73wPomVQTPI9WxmhKkZ6CHrKaoq5UrSzh
3YeIq21fUQ2c+7WIowugnLGwrEsJ8P/hT9NrSQCVxXBtG2vExOlmpf0Ep+sO8G+h
xaSDoZUt+XBZteozOuSH6dCM4wBWYNLD1fOWRvGBjK8QEUtWI1GdWdUVWYUkiJ0U
kHzV/In0ytYZ17xQ4CYOeiFwKGO0wrYx31CJBRGfUDhEPrfx5x5SwbJs8RA6T85d
qMbcZvSVfjvoIL15/+QIP63WhMAkKsQG/MfssEdHoyDhpW4bd5R/h2qFnquxFILg
CxJgOqqKWBRdcKpNsVWtuHzgoTFs2wS6CYsBjm2NdqwpDvLwT9eVkSGk4sItMuEd
9wKldpwNU/0a6gX7/dROrw1HOzjJtOOz9d5P4oprrmeLHK/htbmeasVyS963N1Zf
D4NEBMA7P6OancERpfB6DllULuvtlAeaRcP1H0tyuvB8O2NszVx1rgyhP3Y4Fbqe
RhXar74BfgERAPA289SUPEYBdRXXYTdD9aTAObLHymd+aOUrIBGd9j9Y7pZ0eWXd
8t3WVC4gKlvDgs4sgEUO8rqZsuGsXs2ASvYxWKHS8873AyEJV4jzWQhH/tyE36tK
yypGMwKQVX1p8moAFwVcrqT6rP1Rs5EveVxD+DJPNu9RcAsk9obegSokXUgQFyKV
NPrHHmUj2c6fyjg3N8uiWOaBa42eRc1+ZG7SyaYiHlOwNZiM4EFqJ+qe9opxodwh
DgmzVJjVc9COK9z7KcQPHMNmKglSp3umneAbHvcB8fJzliWVE2HW9iYZO/9dAGDT
5iSxbtbRRpyfjIMFXHfO4L6Ybonm0N7I0ak1FfERGyavEzeQtugPd5eaNbcSP+5R
cdTwc1frTBhUV4aqlCUH5O44UyDT3QFTKgyueUIKW9gyVdxXd2hhGlBWSeCV6iw3
smKXQ6MBIw32a0MqLrbIw1kD1LxaOZ07bKyiB/yZHGdir9rKZXJucGvsXTysHjKK
cp5mWLxkpTtgd2FIhIlf8ElY0PWVHltrILm+uGAa1FOEaMfXfMwK9hqGOFGRTMkc
1zm8w2ncwHXHcarIZa7Za3ImVfTXEJpsxNPOXIvOo4Ugfn1/6vtrA4wkwaEz/83z
Pvg25R43ZtekRwvVxf6RJwffashJqdq8IY1F2y6sPO1u6rZjHUzhxPzd/sO4f9Dn
uit9Ld8ecTua21+8MB+ZzWBSjovlkxwi0pdYo7ccdsyHnMil8oe+WA8cHR/I1/U0
txgCfzBlb8YAIgOstsjuoGOLFz+0d0NiQzuWYIPMe4Y2+n++Mucq9cIQ66E4foJd
+fFsHazLLO3p8v374foCH1A9r0wi5DmP0P3EjoCSP3ORq5bEtVrtgyPxlfzg+UaW
1Z6aMPo8/rN8ZRKB8Ok/sEKDjq6wRxEw3Nzxolb7Wuc2Em4jDLJ/HOvkMxfnaCTI
12e0SWPG7Hirou6nuYtvlaXTuCr+rzNsuiFCx4r8uYjrqNI+BeOu/TJzN0iKr765
ycIH0IOQM18e2q9zVKg5LabAQqJGIB94aK6wRuGQpI0v+fte+tzUoXyba236qXga
Kt5cBV/c0KrJljMYHPv9i57QYGJzylAumL181TtzXm2l90y0Sizzkih6WFBe1cM1
r50lFh9RBTeKKlUU4+cx6PV5anvsKmLqlNngkVh0Nv0G+YkdEDuTG87S/c4cM7YU
3wUox7HK+gX8xg9YU2a/ydk1jCHze/SoOXWVV+EZbrHNBk/xDhTIm94WDwGCkhJb
urn4G9WMIIVhKQ1DNxD6AQVYTcEe5ZcegulA37e825t5Y+spiMivytgZHSCC2ql4
MtomajZqBRbUq7d6ZDaYFxk5sAJCezHsx+PVc1pPQh3w2GbRpf5yp6W9aRcEYfKZ
xFaQtH/pmTbc6Dx+Z8okVuN2B7Kdx/No36RcaVm4tUPvDHD/ygKTbcgEC2HEpX2K
ZdQsffatNFbMnKu465p6Hwc+aGVuApQPQO7ncFaYmeUwr+NoSMYtVMDXbamyqJ2r
5r7X0z9kxj7svwuD+bwYMyAeE6dJjXKQ9rbSjQaJHzGQwdeWHWBwnnN0tqNxbiBl
iq6DFvU2A3w/T6BdoSMY60viOA31MSdsFiHduHPf1OVO/E2KYHNg984Lfept/wPk
Ng8BPm3rERTZBD0COPKYbjke3/4WfIJ0g4lITfdDtbkOH0ZeRllA/ntvBHW9ohMs
VQa+iATLViHcAs0kMWbn31K6M9OadMjwwIV6DYl327EoBIRp4H2NxNHO8gjBERwA
udZfq1BvhM6B6ACi1/Uo1NcsUWuRTAQpSFkGk4lD+II9DmBIjvpcFSsi1edJAc1i
BbNRjia9pcEPK2KkLG725GGEg9RkRx0InEsw4UYt9XGoFcFuhKh08PS+QeZWePlU
4BPRzs+ulcNvRewM3LhgGNOO2ixltoOzjjmzc+wmSPt3fqd3gA89UJCI/VqVgAOf
f2UKNUDNOtfXd2YAMfJmBLa1H8z8a2OEo1VfQKOic+h5c1NPt1knZ78Hszu2Q7sT
ETEek9v24/kmJOrdXTkUlIMzHLVP+5yGez3rS3I4HOaj96YbYuAS3WNryzlyPIlf
+4Jr6mLQL22UsQ2zg2f6mGOknsrJV7U14/Q80Bf3cuybj9yDOVfxmS5rLr98UH+n
2Z3OFtQ9jxHEfYMwQO3EiVT0e2u0M8/rrt1AxX7N0c41t1MlZhufFlhZwSnFIfhL
gAAFYKTVMVFsks2SanLMiJaIGY94b5e31qNKF8vhbODRXaQ9RQwt7IMESBkyXQ8M
eZoiezpJoj1bSPgtvEfpo62PTygZhDIgN26tiXKPGr+Lqzj5hglQcaswLghwDEHL
PfqMOWkDzyZztMyOvaZN6UPtmjUsSIfvrNKbzcyN2KaQASdSCFGFS9NU0O4TrJ2L
dohwbuUcHiFMuwDIlVlufeXrcsB6YfIon1V7O66RL18QVozUi5PDEQOtaIUFjLT9
m4ZBI85Efn6BJImNE8gaUDRtXhpvDbOHtIAtFnUwZUvQ2JoA4pzRAuSZHvfG7JRg
YzfSeIibOWTv0SwLcso/GuKdzbSC85Ay6ukHKdGWdL7h3lM8jLxAy8qu8yp7drgo
2SZlZueJhBL6SriUD3qsx7lYeSTFIXO/jPG8yo9vr/+YgvhgSktSK16l0Hdp5eRF
ieTIAdANB4yE8eX/DIGNMjJUb5Ae6EsJ4DbcEEiluYGU31p6eWb47F+MSDsnPFgn
/9HrUs3j/Xt1IpJ6fTdFqR6e34nBJsGvlg2AZC3EQrctHq2ZLjdg2Dwwjb/PLJpj
z5EcnTVmmoANfoVNBbRwxbRekiaYZ7Mpn+V8iO3rXQEfd9P8xOhz69YKoLsrFrMM
65H74UT/0TYx/8RdHg8lnEgxJeNipqF2Wo+Rl0Hv0hL7MPWXrIN8a5AyJluXpyGY
e25ubJLjsiUdyFts6Gp9pHmXBcMGSUdqDj0FK9BbQqaDo9P7clra/6GHdjaLuQKF
3/EkjFqHG8N6jMlQK21nhRrhClj8xt3ZrKTPI4q9d/re/m6XPaGdvMB3F/UwlO91
e3LMqnoe1gertY2ZVM83hzQcLyGoFxFbAkv5zylsFRi1cLXc4TE2uTt7VL89lhc6
GF7PiS2kDQ3roZSvgoy5BIF2ni9CiMnNEOk6/3ZZofVMj1zNECP3flFuOxfwvdlP
4KN0prZJ6O1HRkXnK63fKRjU+4l61buhWxT1PCI7c7bovVLiSRvF1baKX/v4AA4y
279x7O5/0jFeqTBnZ6y4Cg6H1w6LTSdzukT+uRqkt28GeRS4j/b1dU3ZbnYP6otH
n32vyTTzmuKMwnDZkSv1K+jTwI38KrQvXjQ0aH/+LMLJYol0LfoJv+8q56Px56ow
KITmFlocV23Y73+wwMvHotZDAtRJS6W1Fiqrl+zz780=
`protect end_protected
