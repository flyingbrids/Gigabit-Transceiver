`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Geo/N7fqMQZX5t1M1ukGaVkO71OdWHUjn3dTdqBbUp831aFa7IovCuB8s+w2iqZt
TFSVbBc2YDaesi2IjSHyCsWjjrlXPpbGIwUDR4Nx7++ARW4pO2W/MyPJJlpxNVMA
sP1JQgZAYG9Vy8S4PPpoe20jpJBsmA5sY0N0UZo4ann0vFj430VUxxyfiI+XGxp2
6G2D1TDPlLbBFEEZJ16K2Kbj2BUsF0E42w9gdCaPWP6IB6JHZefCz6S1VTjTcy+9
2g3gDtqhI4uyjyURVE1WOuMMaIH9QsJl0+Dhh73vNcWK3gEFv68nvawadRiv8QdQ
CF0ICRsJLfU58/c5xGGWLQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
WZE7/taDmcPJIEhZkDL/1cqXGXgfy3Tjy7Zt5x5LdLnjudEB6FluTAS4Eu3uSp6L
JaspXN19KUSX1zT6Yw9WTCsoP28pa2YGSwI7JXc+8wMTswoBDO9pwnrJ7/CPsSdX
SAoqxzOGfo6G6nE+DQjIjsH0FY1WhoxindPUyky64XM=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8576 )
`protect data_block
cjdiPoptDKo8cI72p41Ivm99n62G2HJaA8Zh5CUpDt5n3hco9I16BRROqC5lMBON
FGXtIL7GyrJX+v1KvfRxmo+wKpP8iJhHVHnYhK11BgByCusPmUeKQHKvb8Kk83ZF
ocp9QbWwH759UNWxwNywADwz3925Ok0n65PWrlMapk7WFY9Dh3luklBnHcpc07iD
/iVXEO5vf9JgvcL63Xjj0pa2fwrwahRWSkgMxU9xHWee/mlYdXLgu7903vSrwFsT
lnDvTy24j/X50tSWLx42BrxP1YHhSWC4/3ngm5qXGSibdENRYXkB3URokUr9VAmv
ekch01gHMliWIjTQzSZ7rR4lAHBomFfqBoxl5oCbuTPRRREmp7Teprbe5C7rNlYs
+uVyF3ggtt6jGwVFQAvATgIiEIFffY0qvsYXh4L3psawlPHrd1lPYX1th+UI1GnR
LUhlaBwaAt1ABgHhL4Sl6+LmllA7kyAyQXCj1uzVt64lQGtN1Sw0lIRjyq18Ha4O
VjJqZkcoegWn7je7nLhzxFc+jnangoioc1/4a8FhK57ti5T/DejJ9NBOHfociJDM
igKmrcokWGwNwBt9avzfxSaAmOvn9HyVGSLYeelBjrV2ubGVlyi8q2O0qtddR+Ef
+/S4i6DSg24p/StFr+SxsbeSXJ+8nsgMblaDByBXCc5WxV+/qr5AkNb2fgjkSQEF
cWwRjHxHxVtDr/x7qCzDmgIq/1U2izBmmLCff8ktlMnyfXRt+o6WqMOkWRbC9V3N
WScxU1AJ7DRzDvLWlg06Zw8JjWYXrDkRv62J8zTB9m979DXfHT7RJVbBj5fvcdkM
mjziO6R0psj1J5G5i937ycagcPKr+tw/ufJdrigjptVm9FpD+shbU1Uu20LYIWD0
Y03AiLjDisnn+tSKl2tRZJFQ++YuJY9gsX7pj2gEebwkfjiikT9AM2e+C30GFLh2
ul73cyGiJeOypqFEYgL0YPRKA0VNkAwpwDrPZQf4+cDzTQT6DutGCeDC6Ue9zgor
vzguRgadnexYb7p8Ig9/cb/xFZarlSA26LJvdPsTZSYwyvVCnAAsG4vnoIfIHSKd
ZFcPjAOPgMgchnYOpCp/Kh5UT1MqbtAudrdYfKLT2rcqif09L1Ad4yCwSe3fNSvC
BkTacag991Nx0dq+XGDER37/XeuM138rXkZCbrndhy08lMZp5uLwIuBvg4mKhjbO
46JI6/yeKemreofQ5r5OV5Ptlh0EjMWABHZuOzS4MLyt8VmLbG2TEzAmx4VdZc6s
RWpfb8zxXDAvTAbYAqVevoaC9BxxHDHnYajTUCLCLF2rDTJDYyXC9T/eynknVahY
erer0gqtA3u/3UsQ+yBIDlMj/t2VNl7XYiYSbD1DUH/+5HmQ4TlahdBul08eueVz
W1Is6vj0nLoEuQLZW+AqZtXH/L1VqpCCoCyssuSYfbPfgKKoEoaXdTtHQG9MCHYG
N+/PbSoBDPUuNu1PoPdIPbbec4PvpiSloBSOEq5oyc9mmBrzwXoQNY6A2je+7HAe
dFEFTYmoI34yFSIxhLE9qlxQ5iiU7kbLAzSkKehIZflDy1c7QjtJH1NdDq6rB5lr
N3hvlI9sPjvJ5FRXxbTEkxFZZXtFGDs3GA3Lc40bUiwCwZfWr+U5UkBNn+4oouyP
F4Ss+ltAfnKYt7fl7Vt7gnP6ulxrViniIoZG3Mgkg0Di31+unTSN0aP3sWPrZe1u
+Ew6uaMiNHJijMSv6JLOyRnWfU+eLX9pDE65rVyAdgR3NBx5OEEuSAi/axl27OXM
CFUDFDr/GhYK1K3fIEjx6UGlwV+TYea/YimNflGCcg5Ft0z00cefNmnE1oxPdN49
MkQpqUia/xjunyfF3AhHlMToophSYATrIutOcOR/NlS2kWGlmYIAw3SAokxFW7ZP
p4v1MGlc0VImsrS9o8Aa0ETlq0cj9etDtiyo1It+HdBWgXV4XZ9HpewPmZhJQpd6
WZdabB2iCpHhUAYFsMdpkvx91yeAMgCeFx5QReKTMS0yMemiNYeS5jMVZJeyFKH7
x2ltDD4HaSr4SR8k1mNOjs6bL8LiynqvOEmXBxQqH3NkEzMwjEwiI4VjbybJsTNJ
m94m62rmVQv+l3bU2cXima0y4VJSwaxO2rNIBvwSCalO5sLYvNmR4WgPQO+Ivb6F
rXlSUaD2y4sln9Y5Lwnd/3krRWCzSBzGM04bp2nW31Mi8sAKrXdsr6MknteN4rXB
xJ2OOh+JG+xwmOjIjSr90iEH46S1At5NcNsYiEV3JxOSCdhnmymOjhONkb0ttEH1
WKJoe1bKIIHuqMVS0YpzJxxj477RglAXpWly8dUoVmN/CMP6ygBCRAMGv22dX4R4
WPWbx2kMeKqqoVaWf/bV7yFioFBNw+no4sbmRtRr1epWqfG7fYtUUCjJtPbDDq+L
60d60DXSLy6H7rSzEmF24NXrfy7kMA1mqVC/s2CxTCmwd4iNc2tIawOSNoiya9sk
65FDwdvTpNm747aQcBqMgKzjo+8ETmHd8ygq+gJgPBN83bTaHDftKZxiC5Tr3MWo
ym7kfxR46Ku/KateENogNRw6HV9B7GybFHUBuYrUEBM/Fig+S1CfLiyNIjtDXbr1
nXOU70/6/3uZhHuyicy540nICl7ucmSqyRQXPcOpNqlShyMEuWQoJnp0y0i1nxh/
9TpS0KZK/F0M8rSaGRgSwApeeUJPIA+IgAsw3Z/U+/UpPAJFVq3pKanZcEryZHRv
n9YIeIcpNA3yemRJMJrE9h92YtntE/5cALDCi/RB+Hj0E0i1EccHiEzcNVY0gHEp
mc536VbWgqRIziJnQK1l3PSZSpIa3wnwQsNuouTNBJyizyOqaNnBnrTc9G5ziOuu
InhHY45nagx1wNF3atXcScdJn0b4FscF+EMre6XnYP/49d3vdVIxzTN0nKOg++57
TpVuBFEn21Cw6UAwh4WbXgOZNxuZwQt77f+4zd8lHzqa9+NeS182soyWcxpUdCmT
iIi8zc99QllEqvtwLJNL00jjFWU7ApB4eTn6ChHjkkS5OwWXWL9u4afxcN39xyB+
ikiNPyXqVsH1iaeL33C52QlabRRDX5ew5wR72sW9DGT1M4Hc4zN2MmLPj6lelbUl
f6wRAlB3stkdlR9E/sorTestxixBbo6Iot46JrveleSV+fnZzn8rsEgF5C//G71+
DlhEET0sdkFQmNOsgxzffaLTPxjyjn1PzvJIc9lVe73OSfFW24uxwQdtqAbJ2fPd
UC2B+9AyEX3dLyjsaAWNx/tQ81PQKoV3Mv8GFG74Y1J9D9bpH1UUDLYlEr9jJXX1
SHsfsxa9yAjjlno59ZQ9JqBX+2BW/EZlgqd2RH6csEPNEPIFeFXB9HKy1a/4nR1x
qicgEFKGB7ZU9SzjSB9CmzD6ROhgTapk+DvOWrFmQ6udWpC/Fx60/F2OGrg22ReO
dNbSgcRp/EbSiDA5N3h9+RgH/SMvioAk7XNL8Oop5LxpzVeWW1j+gSx9Z4mCOZV5
J86wf+EjZK+5OYVoLDMTbJ33J3uP219Y3yO/ldjYub/FGIPLxcTGm2OhijZvFoSM
mrV2Xb4TVvNN6IEKe1zq3Ydi/CqWL47tWOFJOmjEeWJcoZkk5y9O7d6f0OrbCpCP
3ZzmFOv95Wjn1Dofxv1ePUHeeylot3o/Et4MjdAEURmYriTb7aoz+18/dx8uDfw7
4wTlYZ91znojfv7I+WxiCXCml3/p4UXjJyCn5Yt6D5/QtJTLaqxPUaUlQbzpDnC5
n8qzNBFgWOAYtysLBo1FsF1EYqPr4HimwWxdx6GAGvtQ++m00REQgcNr31L41PCD
fx9ZP7+snPNoGyvImAhI39FV2BA/DHD9OV5KaeKdEG2eqGJtjGS7r5Giz2UG8v2Q
vtQ4QvYAgfWB8frdCtmIC5gk5ceVEsl4fGGO6pINr9LnHicuTR5oulnTpuR8mK/F
3h/IUdLfiluDiWh3ONmFtAQK0i2NMD9cA8aILe5N60LfEkUEVZlBDxyYJR9W5X8Q
XJhMCsXcxYz7sCOlC2giv/4uw6IhNo8YSSl6qrZx0fc2liTUphmrMboMG+ePUtg+
2NGIuKoqDVi5kfUUnNn+bNeOQqF1ZCEr74sqUgkSUDLziAIconno6Xl7bKtkpwaX
UoWYoV4ILbW5csvpvSvewmdozbOAdzZ5gkEVERX91PqeeyVOoozvuLfHnAO1bzAi
M4jTBx1bKviR/m16wItfSBFkIpUBj9DEeD3a9ItNQJ6HhDxo0Lhkze5mKFmtB9rh
7/uJWh05vPvuGufknVfqDydf4s7xFUYfZiwrcEkP8UJVYHY+1st8bPvhg9D/hOPX
Utwh2fsalEGHpjBJygt7wMPr8mo8owA5b14FPbtW1u/VPPrmwqp3t+PvLHmbvkdx
M61RjdoNoDnlSSjTUNuRZ+t7eq+3Pa35s8jKpT6jtev1zdTH2XmXK9QJ3qdE6u6W
Cvqry894gLdXPXSHWmkdrPJAb9kK2TR/BkazRe9OdFhrQy7eKHjSWAJviPfnoJuY
lZevekzRrKeX+9Bfvvo8PAQD2+Myer+okVPmZfXQ//1FNFlUtsgTbfDtC1gJrrJ/
M9+yPAi5NRpZhcwtLg9TEPPlE0usHIx68my0K7q2xsFhP6so7w2lhlhRr/CKG9Gq
hjp0GvEPqfvSSowsQ1lQ2OZwh1S9fRSqzzvS0J3LdRqqvGlGCyB37wRD6bzx0miD
IMOm8tpgA4f19U7e5i0A4IEIoX5qfzgCybBirArlCNBrJJppHt4uuvawRPiJnspb
gTh+QaVOL7d3OMjk/CKdiFbtKXWX4fCnASCXE2ZY7VMbiw0wPrqQhqD4iG7uwaPA
lMQFfx+azH0PIxbs8h8u0XMF8Yw+r2qpbal1TclhQU8IlbAjewsulRbd2d17QIgI
PgjbUthirgJ3s1ZkFz6GKW29Ge/TFv2yFXwr2DpOFYFWREarW5LAHfDFKcVjKtPk
tJM/13jpOWZ+j7+7Iz3O7lLvLF5YVdBUmRYZAX7DZ9QbREix04VI9GI0/N46Kz6E
EA1QyaD9YPqucKW3qQoqLxL3rmpY9X6O85fMHs137WELzVbR3bdcbzzzFWlfAL1Q
18N/fM3fEBCzNqesA4Oc7ykPrEIDr9BUlKWB0WvswsK8fjWgUSGSoXO8qcamQ+Ws
oskKB9awRW6uyKghqvzCZF0+xIf+UcHOy8ajSabomttitFWstF1g5YESEAOqSDZG
SM2u2Gh/wl3raI1DnLZxVqsAUbOiMXJ4oMH9/N5ZFgEBgRx9jPMSuX6Z6i5CKGR0
bebc527aT8Apn5S2z7fk8dTkuHOWq4zETWItZQL2IhhnrRiBjBIbBlxPZ3Uwf1lD
+Oa6SwAgmzSpvvTDZaco8m1n5ebvC2FA7ykl7uvhs5Eih1KFGFHxCdovAGQJPBUo
HY/CTXMQXWe+wHO/wetTEPaWf6EVam06ovK4fWZZT/yquKQo23MoU2vc1g0Wfu53
/cKtinAPS2HvHEPz3SnbMRF+aj20XvXju120ETdrboT5ZNFYka4bIGGiMnm0O+ed
lVixRZyx0SFDC/WOxnDcSX4bChCedAfyLxX4KAiNoAc/O4YIvSoPoVncklj26Jkv
6WSzsAcmM+mzCXwqCQOfXwHFXUyHj/wGqWgZd/N/BH5YhSUV2Qj7YADQ59dhK10e
4mUDKDlzzi6y9bKhJSlEHdZie+779pUr/2xu9FNSESkQ4F7LnYX1fp49hp/AgY46
qEgyF4+2Fcf1kSPHSdZJWaJRzKCgf6maHNKonbF4wV454iFJysZPRtfIvkNXnJ/Z
2tYfUvjGHPHFKKtf/8MeaPka2MaglC+vP0x32WHTm1oukvv3QxUBeO9QBb4B0m6V
dPZEGwGg2i4JZYjx42JgqRSut7vMR1fMl4TQNVHO5uCv3nsgcd/3BMN/E4plA48K
OolwMvrbkGsBWixrl1GFeOasvc1e3iETKm4SHBVm0f1qLfe9Vlnj0GpgNnTDxOTQ
qfXvCLpkEp/uW/DX6C0/c0x3FhzuzIWdsO8nWWBlNQqG4gygWG8HSq1mKl3hVRCj
iCc4sY8tcdXRLM13YKcOx1Hms7JwEmBLaakwfSSBwrlImptapyIbfZI6IVHlCBct
ugrSDk8USEopbgd6cODVhQzlFLj//bcz13/qc1KaaifccxZ8b6jjamp7ZfKc3KFc
1vGFAofo/FZUd07F5o3f4g+tQrYaFeENNXHsCgtHuSqGez41tdBrY0YadN/1n5wX
+EWq8fLFb73AUQYeg2dsAkya8ZbWyoI654VAF7LAUVv99M2moNWjPtpqpfZ/k8ws
gJh3iiSHGBYIeu2fNeBLaKrPaMXRh7fOIkb9Xv0k5cy+EIAGRWGKGWsGWN1Ov9hc
q1llMfrYwKl6Ucd1uc3xweHXSIUDo1uOZo9syHMQUQ9Tk8B059rGRz3BQAhw7zI8
ywhuFGSSE/znmay05c+xideLTB3BHbqYvTOdOSAdzetkCJpRDBIuCPoPnR1yjhWq
5B2qsOgq1m9VrLYmOeDqAniVDpuL+jA/HdXCi6+hAyrfbmAQ00DJlnFBhZgJbBjZ
F0f39+lz/HbWuJz9V1mrYv1kx/9sWvGfGzC6bnjVxbUMFUdGqDjC0J22KLXS/8My
/lEwgLkbkwGy6FyAiJTPj5UNRh5A7AumxncoiNY3t96ROaXY8n7ucpqwvTSbuo0x
I38FeA1TT3GKK017ms+AoXaBbYpY6cWYq4jFsQo8YQKIghrw5bpsSzYxSsW+Rl9B
GIpREt8kaVBsRDCEuXaKwCAZYHRLK2wFGXplOPhBGqiLhX5HqNmjMt3LIB+XtY3W
BCwwc36lr/5iywLLETT0vcYMhSN4TxBiN7gt611FlzLOMzeLNwknpFFMD7oPHYRW
4qJPi3lp8noT3YH5QJEzmSqEww001/RLXyPn7KaXd0cwUPIXY8uPmsT7TzmEFd5j
28HgwWrYD4O4GSHJhN4fcnHo0A80sBxcNWsBXD3PxlUY5+Qs8z2FI4GhFFgcMonn
VoD0K2Tuk/23IbPA11Q513fzrG72ptGYdE/rPDWF7eR8NYJbI1yXardyB4uqE0l5
+xEOllVrhWvFwENyXZUDVboP/I89z9eEEei9q2mI52MjEf4O0p/fSAQQC9nQ6qN5
MPrD9Rg7bV5uLWNcdqHs4i1kMLjOQIDZYS5EZ4hc6vHUfkEJjHTaw4D+BIET72EQ
6LryXwClzsmDQuBpxfh+nf5hxECH0yJLANa0uFugVelioW6id4DhVho4pSaNv4kw
zIiEqgWcbZIbd04867G128HVS5OSadEaJ/vUnkfwaZkO7Rcn+lWkWr0xN1nyXFXd
HlcY9E2zlw1Yv6rDgA+k+cES5Eq0EqLRhiyNHv9l0mVlqq4/ZCzq0eiD6rU6eEYb
Aw+AaLPCGvmo9YqJ6o4mKVVn02qcMc3vktR9vlB/xQZp3fHJmZGf0WM87z+3NL72
hhg9l6+piXZSmurgWsdvfdymxDTwAVMM84XJw5g75KM7H03GF8e+Wh41EnZKJVq8
ZKQTI4b0n8lX0M0piwxNI52Hjve7S5U79Oy+H7gKReMQPFPsw5owaEj+y3OU1hmH
BlmOUGp2q4Es6bBMQ5NDggeIucNv2abclntqGXg5z7ZXMh7hpaCSMGv6Dh9ss7Cr
Am2iuZy3fDge1VdMVGNROCTPzH4V163vES6PgI1eyue48rmhFBULydrvySw0if+X
2ht0wiW4vJk1xrFzANl/L+ZKYeZxBbUJFVqeMrA8OLyYNBwcj9J01a+OOaL/EOrz
TnLrbzIn0MhA1v518qTwJr73SXy1LF6Dtwpvyj2SPOu09gTS3bYfyjuwDRjKQW2u
JURTyyn+64LNAYjLEFFh0rNAZMfHQhR6UYHVtT0TwcKj5A6C7GP3NeOJhVBPxPkL
8qg4Q4klzIg9AM2vFXswjW8DPUEQYibVeCM1gr1T5ymgz7ZK7McmLLoNgMEirKVm
54lVfzcGG+L2OQt0Yf2/ftvYrVdbvb2sZqvBKUNob4gGQ6SbzYkZo+12s9qrI90K
aQFmqYIxDCoyAZAMUUH6PTPSWVS6NkhyoHeLTToIlx+OF20IMTE0X4IYbha/LBkA
ZHhj13cY/RzkjrHmqYLTGv6gZT5EFj75+fY5aPD9jBGVEhfXxe+evMZTSWSJd4DO
t7Wa4OGsZvp4SwJLauSuOZdab2bvS8/qVrwxVe72peGX9goTkdSZwKChvFwAabk1
fIRCBPWReWu1CTRUkTkxYrlla3eXHIJhWhkvmr6p0UOQ1321FsswMTXb70nRHFli
gwkmeeobG6KoFsJG1P6yFSFbzSEclJk3/ENIhrbJoObhVNgrJi/F5WGG7FDqO+Ne
YmBJ8tG6icBXCgbp6ikh9cyxyGmQOCJH53bhRcW562+i18xIUuuXwaLFm/aII6xd
eDnOd4GNaTl2pEYXMU1JPlwTOI4pZtI479pTRgzCPk+6rOQrA//JItNgVJiI1FvX
re2tN42LoSOFty6r9RcdxRgGYsvwNYkoEcmT7E8aDfelUNmfeiHhF0RdAqUtgAG0
OG2y5HEWJPpgM6Vr0sQqd4rQq7QWy++C92RwOEGRmE402DIKrfhxEMishhIxLd1w
YWCOhhAkLWhxwDmObP9GJU5y0q/RtkqEcY9BLMP8+r56mAP2D8I0dtRn+OLOJbsC
YHpkgOaWxs+QaVO9XDp4yq52iksudCOuTSSRDfbKAtpCxhdQYWSIMu7muWo7kZ8x
4tg2KjPmgQtwwxAZ+9EGSUrrCVLI7xfsmC9ptj3/YG6QePJ10FW67lmz7oxLqFJ8
rzEFhFi/9YX2oF3dnhIriNt+sE9c+gpI+K7u52iKjP2IBzDe5E+9A6PMtf2dyhXv
8bN9rodSUnC15ko8Pff3+gEzgOdRbKFbppWWxAj+95r/Ng4w4eeK05qe2f1V7F0S
dU/pr+3cuqCvOWEqyTym/j6DJTU0obxNFiuUKeJ9outbSLu2M/vk04tTFrFs+YYw
Ue0jf5Z1WsLZTxj6CJCxSX98LVh5agwLBlJadKe9b/xydxs2oYQJDv+76hby1Azo
DhTEa5nRAd893xu8avnGhSW7/q1UhlvrbLySEmASxCuCi+DbeVDvode+DVuLu/2n
rWETFKIprh3Nfw5qs2VnjE4DLG87ojoy8dJerYBvR8HrM4hvt3tl/R0t8XzYgiuT
LLhD0RsJnYEWZ5uOYT38Owd08iqHI7b6UZD0yH0EsmO8p3vYrSemnUbf5AU6NUKW
u8oRy8NQeciDuAT6mPEL+dROA6+AAyRRHwqVWGHUcwNlbGm707LdH1PFd4zI/vF3
/U9msbS1qiJj649Lj7qI5nXe/xWG6Ulz2DtDb2tqaopmq1tz9OfBjnHG01MCvvaY
4QD2+G/6cPx3sa8PPonc/7WCBfs3aqJV2lnXFZKrLiC6qMyG3EHSyw8HHu6fkMvf
gWR3mSr27fi8lns8xzNvPwZmA7aorjOcYXxpgcEDioAkD0smTm0vW4nqkJjzlE5j
1Svg1s4+SuXsezjqn/V518ai0dhT/qd6K4JbFUnUQSPn3J8BDrY5W/F1CR19f+NX
5/SmtIUyFVIMuWaDAk8Od5Zzn4jAnbq86G3EY7DKbT7wGrkfK6/bvS0aU2s9FPRI
PvXq//jmErzxBsDo4+P5czXdLhdiWpyrHi79KM4h3hQbI7PIP0umDMbMI2zV4eqN
vkM5UcQETW7q8WJ3Dyu5xR2LGXr7Ve7c1yN/stqnNbJQyPbIGL0iEcyNh5vlyUH8
i8k/Wafdtd6Yi948GJgkCNSaL5nIEBxzFWqmVHWVRJPSmLZn+2J220fKEm49l/qw
ig1bpBY9kFxvua6dbAS703bngwSrz4x/kIcaPzQmwGjmNkEMo6nDYh/Tpr25dNlW
Mjfe9WMyCo5Aer7ZaG2r4HTgY4PQRGzd4+jNmJoVZ+Gfyulk3krNc/HR5OoFOhla
8f4kqK01pSpuMiVBUHHtLZZOdB19v9qciABQ7CBxdyliMyOZEuB3ZKokl7UqSZXv
BOXG0/GUvrTlt1z2Fu9MNGugv5BNKwr+Js9yeVBFUbNgVyhJNqrLc5XBxY74u+Is
+XmZw0r5PkrzUtP86gDHdewbNpXTWituOWEF026PTCsSjP0SSf1Jm9Q/7xUySJzQ
0lJDabmjLCQ3oQkwCvX0JLSalU2B8y1PXRaMN23YQHOGQ/fGuoTx72cHCSOt6JMT
7qM2jLJVUMCkg4V/bOIr0fjDgRYCJeYG91yQj2vLhgoxmRYq+2b+Tmu6UP16PWq7
nYq5xTu1sHqwz2eU8gGah4MFO2FbSVhWEPy+xj8syttjA5JLqbvPXGDwRUFboeud
cePe7EjYcglahrYzhpiJXSm5/dKhw+dMfR09zC0PiBjfF32ImcnRyjCcdAqUhZT+
pw5KbJcqhCntug3Pn+HJPBFo5Z5bRUOTpXFPKgjBMKFHo5kbinDxJmt2QQIJd1UN
PGQ7+pFKz6s970/qIQIyudv2Zy3FuuF8WDwtNKvfA8EAANK3Jp0j7moyWtwZ6qnm
aXAVL1pRSMi6GJHhYEUpZFKz6Jckzsu2tmv9G+e0oaNQ9c1H1wltSBQAB7fTdTQZ
88noZTqv0Hm3x4D9hZjvasRY3bZCLmINhFVj1qRrQvc7YBzt4R/BqzHtWu1lpula
0XAFIAUwXX9r84VpRI0/LyhwbV/tDLdhFZmIfkwMDzxZVP1arkq4ZM1xE9fkY3X7
/+MSdkekpNjr7yb2O9x9S37u6CxW+1zCLBIAVoE+Hs8dDm+WhKJxOzh9MmTE2qBI
kUZGy7jv/Q5wDol8dX9uWRHtBaNXd7NsU4jhOWnm/5TVYFXV1pRlAkdjXG3n7ldm
og0Fmab+E8tGH1/pP7cpioRAK92sQghnJcv0gCNU9bi1JaVxxtvK3u/g6sW6JcEK
kEFyuYp6mlxc2dQs4WjPjCaK/NLCfiUI6jxZyN7fEZX1cAZyfRRWA7tXidmkvgtR
xZZt95nAQBEtQuKo6P68aP2jIafuEZ2z52jPLTI/kelHfYEt1neM26NCqT3S9hel
+PSK2bzfC4er91iJkIbhS+Tvl13+sLcW5jStmJVuQY4Ja+jCRhSpfTr4LKMHJp3f
qD++qCNFUfvv439knKZ5wMaK8tRvTCUwvN+lODo0CdpFwKkAz1TCplxXEEci8NDT
KxuOnq8jdYoRYEb1ZOiVy5Q6bLvqUF5p4SdQKrEosIhtZEUWpbsinParUuMVRlqF
vvqo1E1kGl4rIqwJLbFvNaTBLXeTr+hUEZxIwqkt/u9vcfpyVBByVrXGLKNwTUgi
9AhMZQjbWsgCCYiAlV2NlTqDbJwAYXfx+QHy7UHqKHGmyVtFPaNHClcwBS5Wni4h
n4fzIS44oRQyXF5y6DQzb/G93UFqJdbbc9FHDu/72ks=
`protect end_protected
