`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ccqusA4EwxjuziK3Tmy6D4nQ4aYTiKzgZ4foxs37du3pJKfArr0tCzkK3Z8sRVXa
BkSJzeckC9+Ts2jsXi2ybuEkgbWR2eVJl6CZEnXn+YXnEMp4YRzDM7yrZ2IrxcQU
DVBVQgx9sdPM9LQSgX3l2UcrO7dYlr5i2aYY4JQvcFaqxQkLivJPfvgvBYEFvPa4
AKB4OfO6LT8OgQWCugpM8BUKeoTWagxQDR/lUFyJWjp/aRs50j/uzRpavZqFy3dv
dvzlB27gf7aKfvWeBq5601/lxLGzvEjnBjKGsM/SfbOrHp55/5B6v7iO2JfeSNh3
zYuYFVelBoOkBbyTbnOm9g==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dSs20KYGwufxUCmRyzHR3Tzubm+lhwkLTU6hTjx3pGjn3j8FLHpQOlybAo8o7jwV
entFQT9pJf7aMu132Kemcz7SRFBf2illDZfJprPNyQOZ3ZWFB+iwYyi5ZeaICTvp
sDQ/HlnMvumXDPiT11OUXJ873RfqBvQXg5ezNuY8wwQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 24256 )
`protect data_block
1WOLYEBHp/SCoHkuNA3I31piYQexc4754QF5gOk2VSGmv9B1xD1UUHoufvgbLCd2
DLHTflDUUWOWLlySjX44aZXh4mnDwBW7CrQ0MVPyxqha5+6XGZMTKr+DyIf0628F
dCOUvtyyu6WAyQ2nzratyelhSmX3P9YhdZ6b3On5LnJfQOuimCyLewiqz5Nol+CN
JCRX13LcEeFnIw38mG/0dqqGghm+hHjjNg/TjcBs56/S+t6GKcHiIW+mQrWr+3Rq
CdXs2gkDJ7qgEBqz3dz0YnyLOyCMMW15GZp3HB1dlUDq/0zuutefH1sRSQrPknFs
bcvgzL7gSQBwqDpBCqWWKfqwzZJuseHKrdtFoe2bjZEO1Twhimv1jFBskbFOjwVI
mENCrNajjmJA2ZLDaXDKfUnxbePfgwKGVmZV0EQJ5Bs4qgSZBl9/ZmnLsVXIF8FY
qCaZni1Dun+suntFdYP5+hfTOI4Cja7IUEOlSEBApUJoyVo0tisYbQOyAxS6E8QX
EMQXKZ3j/BhuNDQi4lV4sP2IEuwehm1C49+E7KsfjcXIHkHdK2fmGyhWgraAg02S
7uGoGIej0UcYee36oH8BAyyUhTmnew3ohOh6/VZ+VYnGm3KOyLnpIc40tJiGyK7U
N7nIv/m6ugoubdClFX5LmhpRawWwkeuCdyQxUzPTe+iEbIHNl/o4G/Eyk/ckp0EM
Zgu72YUtNiTysRTqppbNxQ5Mcw0gKsuJRNMztNgPntSkc2Y1v8sLQ8VJJG2YNcb3
G5ZNXQT9e4Nl1bp3YtUCAVLgCf7hyl8pieRN9ACqdMcR60mMqNgB5WpoOlfFdqwg
etk3pDmoM2R/tI9xdMjpILayySFo6Gb8GQRX3l44X+EmBFrkgOKvY1AmNpEwaTuW
mBtJ6xXYEke+QNPjaJNh3wCZ6DnhxFJ0JQTskgDZBmh+DaR24IRSo8a87bUG99oy
yoSDiGjfNSMiKQAXHpBrpkfrQMDRpNqMLmDhMTyVI8PwUWvpufhsuBNLccw/UvnO
86eaB7UWgbfgqLgndMF573ajQK7hZU48MFdU9AoTcrCR/sx37ZaFBPTsIca+HdqI
AFTTy7kTqlHTAv23f8T/PNOqS+Z41zDigtRue4mg5IjBbZQrliHgHHOZbSnrWqGs
24XEpBnxgxZwjj2zN4SbnOKhlbc/OnGZ5VaIPt95BK953Fl4JWbxWdcmim0RG4UH
SuaduOUSnj1ExAoQukT+M3B5MUs8nQfFnIwnNYNQczXPbOeJ1Q6TDAi44r7Pad7l
RfaWx7Ki9TzTEXKBQD1OC+8fn92W72w5y4fkyIJ2/DWBVbxQ5rUZHF1t1/JEzf2J
5yxADbLpuUUAsPtwY1pw5qczU8vmBuGSlmEtcZhhW7pVYkTR2H7pNkh+ExVzsvOh
pulWdv7VODqsc9UDLXeu8gCUSBjiS5o4FoTzlig8WuVJQ4r6lw/PphkKHMmdkVd3
x+6D162RYJfrM6dabxFyVM0Xro7i9idaGDzqK6nS8re/2YsHWyPBIneHHnttE8eC
d6Qeih9KIK03VIoULEI1Hp/KgF0XH46oeeDoEeOnpadkzvKtZzk/OZegsnD9NOe8
nMBShG6XMWDeK9ebv/OpPemKk+PkmVa1qOHhAGSyJ2yb1Pkadq/Gv1QsTcvII8cC
USvkC/Z256luI5JMGssGy//88BW164whCeBqdH+mJ228hm4mkwfIK4kHVPs9Sw6G
S/XRLNL1WJYOmycTxKWRuUPt0ndzbEUwYjRX8N0sTFB9wJ6OzIhav3P5Q+JgHSJe
3fOe6Aaoz06u942rMEZ/0ISJrKRZyLBBCAacwkzZAuVSaAJHuFBsaz+DFPA1xW63
u42WbgTB36vHqMNZWsz7y6lo9sK6iuagWmV2w1UhsfMI36llFDLW0pcNrn7ni4Hc
Z4hx0LHauq3SeEt7XZ1X6IFmEpqm6Sa6y8iV350CrpxKvymGCuAgd7SSwTwBd5Qm
2VYdxQgjCNNEQ2A30nrB3/MNXFVhTZIsS7esZtlbgYrG8bCZIH6DikSQ4WlRI2h+
9xvuUjICz9ws8qdwrW1/lu2OnyWBKf7G/bJfXcy4rnlGcuN9JNn8W5zujOTRcgIu
GrIWQ7OYTcY+6eCEQ+3Zxokn7PCznKJyFkMRQ2m02RuHr2SblEjKe01HF2imOWHY
Lm2CrUzaPMl83iMN6W22V49r/72AL83xh2IjRNoa5fZbpWPl9SS25DmsDFBhMq7l
kMGr4RKkXtg5Mw+7GJS0j1KpoGRHZm7mvWVZ2rRZbR+/LG5I6yuhEBDlb1Jzsa0a
y8D+/RRzt2Jynq9FSNekF1yLViADK/TznR8rEn65QiYGbsOOKh+/a1Iv5LtLLWFc
pmB57UyuK9rQ+/gzJIaVjLj3hUY6EeNi5JmzkFOjC+lWtlV/dBZ3Uv5PVYKMd6fj
+yfqUN5CtpHJmHm71Ae+jIc3qF27Tb39zDX/Q/wPdI5YRDyMFRVhCTpPuvSMlMoK
pP3+QZnRS4teYg4t6C9JlvHQ/UuU9q+CDwBq+8UnymmBYbV2U7YzTUbcP1+MXPvw
m4nTFkQ1itKNyRvUJ3qaGCOBJH0BC9mOGDi4o/nAXIWGS6rS4GqzGuXO5XVExAKy
24oe88QvjAcpwdFecHjL9mbfoAxWY2SJ/lqb3W87sEfIpN8aAMvt1WsIP7NiyC2Y
w5UG3V9iiZlWLoBVcabdJ+mb33BrbnMpjsaCQ2CBEwBnDEL6/1eCq7TciTFxQr3E
NiS5TxJgvhgDNCRWmJrhW7VGK81z36UPXd+/1ZBnn8kiIF7ET5Oo+LBpdWrlM89T
M6FxqTfkk4ClhdMkqrT2ZRyQlbSYJLmR7f2p7OaympmGpUiVx4IDLNqASlfVpeGv
73LywgsIvkTXx9EFwO2NWlo+OwZG4gTpQXEJV0NqnUf7ds9okN5gUZ6spnL3IZVy
KyNcYZB8LxbaePYa+wjE7RoqQgnaNZXE85eTKyyb091kH612IdahkJ81fiQDISCU
yEqWIJx0FKZHAu19fOKZO6Y4VWkO88EViNLb68qRsE9ZxTstbpS7Y2EYkvap1IU4
uHOQNk/IFt5h1X7uyWexehBiynff/vKoQspR1qHUUWfAOJtK1KGDbDInpL41BOci
OC86fZXYyN0xGGqrbyypRuX99XmYeoEEb4HBgzVAOCA1NU/M32egtbul1fJJ/wws
/8nef2u08aYrdrEyxgfyo8VTAOaV2QD6RdfcJ60MjgoYxHRnGD9sOB5ky1Mg6kST
GmFL/NAWeVLfQYAHocCfiC8N+nr64ciBXYGEAsXpBUKXNWchQSizgpGDEzDTJ6Le
Vr4ta+H9X1Ud4ShoV1bNHSTJO6xUSrn7Cx/mCSIldFTFC+gFqAIBS3k+33pFu9Hw
tXd5iLvypZs7k61vP195YnVBZ4ra9kY6ibdp/8Bj3cPLxi9jkfUo12LvjoAALLQl
Gj216qWohRVp+Ag5yotiba7xFNBmeqLBDYf5Eo7qeWhC4NAhgiGxh3kzUuZFn8ot
VHCxL+ktZ0cusyde6ZBuh/OtgrtR62A3DN8WbDRCqkIbSWJKr5xoGh+WvMzemGJ+
gIkW6rrr7Pw225tF6IMT5L/gnCJdUvHVxsD/pHARQFmCZHKLobOfMTYP8Fsyg6qS
/jW6isQE82SY3iAcP9q9NchKvuJ4Dpof+FIEDrprircvQqSskfteDE/L2UsXyIhm
LvytTosBL6u0uJSOtSIRHEpZWOeyUB7X35/LtwaaayolOrX+1SAQ8UFTezm5B7Op
qMt3hGsHogOY6TJpaLUlmJ2JwzN3r6lp7X8tmMgDoV9oXzJuXMO695cpwoYtL9tN
m3M3H54w1wRDMK/iJ88vzNrgdd+qvj7Tx8H7Xzdvc2sg42rCdOkm2c7DpKv3gVjr
nwhHc+p8cEV8uVhUzpgLXx33u/ogK29lY/T06Jl67WAhFcqklWJ5fWFdSgYHOHuU
FAEUDwpCufXdF2DJWgNVDKsbdaFTIX9zbhC45zt/hNA48dJtHuBQtHPeROXZWsty
7VW/BCSrOzjsO+5fNvhlEiSsVMtIua5HkKqLUWzaDWOqH2yu2ABKaGgdJeqX4Adw
0I1CKDtm7Q71V9QrE31cN0ehUSt4w8X2NZ3X3Jb/gUWUeT/VTja5Q+T9S0Q6+Z4f
vX8ZY6IQSTfeeRXKAQOHVYeMeuMN737GN1MP79dkK7ichu3gVjYQBGi27i3leygn
UKimVaFJHloTNEXWeYF0qd0zdZokAmHm/SSSZasBXWikvrj/8EF0AQ7l56auh0lC
Zq/wK0lh5ZDQUD/6BaoyDb89N8dpzu+ZA9FK/LNlLnY/YMHv8ZImWz7bwEZrsA5U
kvyq8Ts8PoxUSAujXP1S1rOeUazSrYDX697xg3FuGHa+SkEFgWOlPeD+ApExcFoE
AW4Wb41TkOWCmTbsdHXjMJzpB+ylc9SjhhYxGKZomX+oP21MWa026P5IyYcUv1QL
5E/RxZxI450v8JVtfEHgYbmuK3SgTW8+jnfABeFK3+4F63t9sA4YuBgtMkDiGaM/
5MOdA5RSwYSQQKOa7M7AW43RPWuM14vf2zbT3OEM6r4wvXhUdBpnTCQ6UdlaZ11Z
eXKhnGs4vVW+Eqp6CmJLZ3aZbCJb9FrylzOkqnjs4Q8ZXUl5triobEQAX9yiBHix
+sPHnx/M2PbJhWd4OS0RQIYsVzbQZww5TH6WRTAj/zsCAK1oyAwaqDooUA2+7La2
IZ8fmYeER5WBW3T6Hco7PnIkd0AcUs4sEk3ka0M9f5+Wa+492xhZzvS1h2GOQPE7
qtSVFRuwNUD+PRj4lK1jD6olZfL1Btrx/bhsifGYuWeoizoLfxaonx83Afyo13oN
bP89kqjYB2CpPAdZHCc9c0rhm5aLZHz4M1AqxyvI46MbYD+2KHEC7hKjlRVVYDjM
8Godr7qs+stUy0aBMkb6h39KkB8AR4ciJLOMzjHriKuLsrrmiAQFjk1m06PGHoaA
+zeCWixfZblKSzR+MemPelfJzfflQyUei5cbkruwRPEYPZliPq0FqUgfeQz7t2tB
KAeNBdA/e8h7zRRQ8eChBI3SXp081LgQYqcEdYLb5js+x5/MJjbDcjlAwCG1Z1/L
t79tUULWk6XVsSSk10oVmXFYuWsdNmEtCDd0Pclifz6R/Mt7bkydkqSSVTK36JT9
3tuJUAb5ZLq0YTC4UuyE0oVpcML7qvtQJdlRojmFtkXgY3P9dLVaBVCoAA2ZTU5A
kMpgSjM6stNJoRKVKy/08y2dF/2KlHGZMBI/5Sg4zDRJDzH8y4fhEbXaHLWuoyg3
noDTJaUgv3YoLBROUtQiRqjtbF3LbVr72K10gkDcpcgXJGDRGAa7QOXPqY1Uqcpa
ztVimyCU+JvN2gfNc23vBAr6FUsUdx80sT0cAKntnpvP0G3ahcwmFe2Bnnqj67WF
ayCpiYikSpPsmVHOPnFURkDBzHSY14efXojin8bHFml/ccFsni3N3MOQqugMDYED
Y1jNTwWbO53SEkC+Swyszf0r4POkM48URV+3+NIGkPVvlsJiSU6ztxqFmgRHfuZ7
TYJIinEGDJG3LMf3iFy0Zb76ArMWNFfGiGo52X4Nd6Qw5K5lPtGTOElcWA6yNYjp
wAqX/pi/1rC/km96iAyj5SCR35PDKMjxbnoyvO+ZRHyHrCSKQmVMjrXxo3oaxOjo
g8cr4IZuPxDeEnLXQbSjta+MxuszdsVXPZMw+qmxJsHz9reKg9pgAMblm6Qq1fM4
kYz15r1vNAVqKF+5f7K4Ke5LFWpeL5fJT2PMSV4XmXrervSvsSCenW2F8MJyDZh9
HuQmgeqUx04/qZmRruW9YabeiB0/2o0Wbw4JCNhD2Im/fWz7V8XmT3Pza77++P8a
dg0gW+1WnZqXU/yuA8DP2kLOuBIbfmX85Yuo73vcdww5E9t4/Y6/C6YRSJTCFylJ
36gKThxd25tUs8kojgnwOrDVfYfR5CrDQZ7DU03JXY2Lir7gANa8SQD4lwWKRhH6
vFC7F1QvUS6N5CjqfkGFeVG0w+2SMTMD0mVez3P4DLyjmGBLQddSSk5dm2Z3IEmG
kXP7fonAB7nyKacsZ8c50Wvp7QEsxYfMMLNU/PWWGGNzGg7YBzvr468IxwGwbH73
NPsjCOzMJZhw5uS2WJj+gdNFczlgHeVVBWXnykVpYH1v/3h6vMJVlTCbmmLl2ryi
94EvsQ8YCfmYnkjbhEK3jlpHrp104WyANf76niyTF+4X9n0EB3A27WmvFAW9rWgL
StXCO2vAkdenr5IyKBdyX6y86Du/7Kf9fWlfovHDVLSIFX8FaWiBVK8twmhi+UQG
thZyppM4EAMuH2v4v5UlN176S5rd+kHkK2m3U3piwbUUP+NUgdBnq7+lPX0xhidO
208zWoOv9IsDVDbQSjAVPzvXXmNcOemPLI+9Scp333vgHaVlaX2NY/uyiMBWrX1s
isaT5knoFiVMyK/NXAbN8oPF+DFGUjBAFu4B+xbyt3+GWtXrC8dyMOv+JoA49L38
g0Ku/mZlJgv4HmPOLMEyTBrLffZtQtQjWv/8oypPAd2e2vE2WbVRK1dQx8TYSKpa
pkX2FgAfIbGlhcwRtWIj/6MBMNw4lOldm+ylCDjc/GQE4BTRpWW9olxHEic9t9ws
xrBKubR9OUHbPC8y513M3WsJ2IoMz/pwTxXzYLZahzLhQlpVcoLX/Y7vEcHYbzas
wYtUtFwj91X4/kpN2FcNO5VO+LwYmYtPcN3TDcHAXS9YZHthBLsaBBhjZThy+06g
E/O1k9Cx8qiKZC/tMZp3hoMora7dyGcbrWEs/NRc2z7JYS8x60e+XkcHNn7WYSCT
dGNW+fkjK7Gyi+HjrrDkLJNJWIVEilaRp25baIF3FCLsUup6ebOvDLIUNnFNWjOC
L+STYAEaodjhW05HfD1tKxl1AKAUJs4V2XddhSWZeb5qsRS014OGXpn8YFFVdv6a
/ynq82z0XMWKz4dC8KWo9Y6qV83dCsNNyR0hMzAYAvCMtge0shCMEPPeg4H39y3v
BCl4qWvQzbByJY+Ntfr/qe61GW7/BNlL8/ZbAKUhmfwl+YoCgE1RO+0e146rIOfm
qGAKXavvIj9mAytpnGFfWBhxej9t12HpMEH+jc+AUwT1fcJbaHQf3RzPbJ5a8WtM
6kAuFr0tFnGzApc7MlhioZrvJ/F7hSIE67sSPepqu5Y8EimJZFk0n7sOb5+qiUMp
uLIV4FB8Rvr9Ojqr26P9qxxJT3hiilbgu8sp5s3W9gsb1Yh8sfOKRZ1KkHFaYHyT
E3OGyFnzr9Po96Y/VjHwzo7CgZ0PdJ5gdyS3pz1tAv+OKhtfp13CthcRuyIEvs5w
AjMpgScHGPXkPFCXfenip4v/FERVS8sse7a7ThlJn8zOxdMVuKgrQywR760dQtw3
aY1lvsVUKzudvaNW5Xg/4WjAc6hqRUfRqGCyl2gS29niS1Lz2kPdCHWU5cYsufl0
Qaa7NFFpneoK8heMuKCivczC1XrNONAIsRPX58uFIkJ0BCSjre9XPwFrQGS2AAUT
8M04ef3d3Abe6Alm1ePzTE7rvSxAf4IK8sxb1l2uB6oMa63Z/couKuGu5qRHoHlA
CpaAI6ahPxohJLyGOcwgBhcrjKQfX3dYELze+5r0oCFQUk3HjATlF8AQx7rz0P1j
DiW9lsvB9KUC+aa8hXm5fiJHBsb8pmozBuDqkE9VQAX6v7xAr+Ew3eSgWZ6ihoyo
Uzvgpg4b5CDKEp+U7jlqUaCzizaV3zagTJzRmnVwofsXHUYGeUQeJMMmNWV6EvWp
BIDfKS8fkcl8IyFeaQqYSIFy32eR617zOqjxquI1mLfVLmvHK2+Ry5wEt9v3PkY+
FB4bwqd/c7PaSnJNAzL+rCatdlloZqJXjuefyUl/o18J3DzA0A4QLb73H5Z1tdaA
HxyWzslaIO8Pa4Io1cmbGX0HZSOAFwpNn8SYHl0hqY3fP38wVTL357pq46WDfmec
sdO5Eo1KHpgMJZ37DAdJ4liBXYQiXoFlwoWKXUL08Rpj3fgG2yuDBgSOyspjNBfd
3wg8yAW35SsQLHrWuSDuonrlyAincP5LQxxVuphg3nhcQn6oz9CDXm45br9w8KW5
fIT9vuVirFofrjxOGCr5rGSt4vN7Dxz7h8FqnFGYnRCtdsZo3R5Oy1bHTgIChuAF
WcZOMM2FkGhRMfcT63fdQhH4T8zzidPKAB6W9iq09i1Z74G0Zlvz1ZqG2f8nlKMZ
SzebXzvzHwja7y2e2PzJ0MZBTY9pSySUNRC6sQtil2Yuey3PI6m00TtnxlGipJqk
GiOyML28W1qv4MOERLoxDpogyD800GZeFaSJEuLb7ZsZ4bj388xOXiMu2IGPE0hu
U/mcy7kfj/0Uee2DImNEJJ0z+Tt3QZvey1/2YucFbG8BPUDwT4BPQ/uy3TUeloTU
ie9oXHCWQKNBC6MMcU/sW994vm5Zv5W8o7+kBcTbpnvjgvH9uFaE0M8rwDc6IfmZ
oDOM/3VBir79cMWxdug9MJAwdtWdQeYsfOYcmhi3nIkOaRiluTTd6a7tntH102kE
5GmdPmvKPfjoJ5E5aHdpxTRQtEdG0Hg3mwyNeqIeqDEZdiruZjOQJtJHXLelPuHo
tyqlrprfDh/4Hk4rrMu4WBYvqmi3+iP7h/S/aEWIpI03Nwjfkz29ZrR2xYySyB7C
WUJOCFQIJoTLNAFalqd4kBNC6tuiP9LayJWPZwbMYvS/MR/mkD5S/1Xaw4xD7AsW
p3uuxUPUomfhmTxI7chTmlqcuOUYbvanpzyV4s/mQbAz2J/YhRgVZoU1qf7/Gv/I
M2Yr8G5TsvM7GnL9ATbaJDEKxHwZ+oHYuxXgMbhMrjYddlUOwG1PvHA44YAt2RWi
jRpAMLXxcvLZNZfmzNjr373EHEwXwdCzdTS0HVn57M5BghJobaiIp9AhD5wr/e51
cCD4cQ2XMCjmtwxZEtwuPMnGCWEy2SKidG0JyOQQm1fVxqI2Knt18X4pdmfXk6Oy
HQKpgv49C+YCJ/halRs3JFdJpEEx01C197liLyFAmn/zGNE8q/InI4v03NFGeRlk
t3sHJyCyVujQjiFB2Po5SMeZmZk0iFnKNzXqDb1gUm+RN0jdL2efmW2Q5JCaknpe
HRbntp2fFWQZ6VeZJhnCZHq/ZUK+Chs1mnhOGJ5tyRElGcSpoyHE5qCUk8YPVd7t
Mds64Czw54p62vZ7VikMggkHYCeZuRHa+xgpzRulkut9vJQpR70tuD4IPYk4i6p8
Dr72mmI2eI2X4UNc51wtls850519IzLTfY9G5Nu2dPL7zADSFOCrqrYRA5YByCQF
UIVKMZe7DEz+NV1xO8nxVN1NyYVh1JCWHivF2+hilf9q4mfX+/fr61KBuRADN1ZF
whZnsMa5bVE2yujgtFrwwRJlJ9ISX8V1pMmmbe/l3TI/oYByvqwVKq31XEl2ohJx
YY86MA1LCFrHo8+lx1GwHz+ClAIAKzyEUJgb9+jqYW3Fu9luzm+6PN2krM14FEPi
GDE0nerqScLvKqBlGGWxgKZGwJHWJFz7r4Qj1msYD41VxfCWNGcrnwkBKtX8cfEk
Ek/BNSv+qQRf00HwzQKDveBAaXZcCOFVQgWGyRFfbBseOxOjlgXmgjmTjnNXR0fB
Ve7DePYwAuZyyP31iDaFKZXsvIRrMMq5RILjlBM1tO+t/AS8sk0KDtfdTkX0dKfd
7VfP/LKOpzyUOczrcJvM/mYwTPPxhsYq++636usK+ROA10HmnTf0Spggqzern9Fj
3/K6sMktKIRiJX+V6Kahlqujkeqskca+j0ssZLxPDtNetXGx14IegFuwNSqbEnCM
NbZ31NZU96ZQq3pOfwlBVSBkv9PWg1Ux+b1JhZJoR6ydvy2RQ8AfDF010PoV5kdH
6ZEW88H4nd4dgqb6Sq97e5ybVD7lIyf8RaWDh34L3C0Lgf9a8qfeNby9nE1C9iAM
0UL9PCSPMSf7i/Ze9PqMFNrEPvqO0Gok53lYmUpjWPs1sXDGeevj86AmQNGFrVeq
UKszrioA8Q/51JrOJYjFzCatWQXDQbB8dXxLC5czjbf5zl2P6kaWiFYDEfS94zXH
HYb3BXCmXi6NJ06kUzdEcQHCCb0ACnGAzG6nR6yK4FYOr5wg4C63APbYw0D+K2GI
VoTbLN667YmHCFKa/5JO+KnfEXbf8na0FF1kCJ5ea7xFSy2p4qsnagE/h1VzoKpG
DVdAsTTTBctEYoVBZA2dGB/F4dgTK8bz0IOJUvXx5iw7oCq5TnkiRYGxTIf3zcoT
20N0lf4/FbqHEbM0wdPlUz2dlT5Qt1maYtF1L3Tv9ezZJ9L0AaNKuuwMaaUJIuBn
ROLtFaHbrqITP0A0U9m+BVfnjOd7Xh+R0hgZKZXqt9VxOsn5PN0eykj9hHwzEaH7
hJNsZZgKxi3bHN0MvVuQ9tgVRcXCNdlrVH5+p6rhjFZsIwWmzXFvdoe/ShWU0Kte
vw3TT2b/BBhgMoWMZmST/qe+7SPFzBI9vSzRBE3wmjsVoMki38lKRH2pbAZQFd9J
MKd10Avsn4t6q4NxpVRwAKIqP+7r9EX7wCZu4mMy6a6IT0qOlcLdT1sLSnQzfmYu
ACfFvwAzn+MMJgB43Lk3aLUmLQ5O1YjbTIBZQ1DWMi8uvZPd+3LSE49uT1oxZaXf
bAdSZISvg2peJ2kbuizuE4/Q9GNUSjnwtz/KbRwHz3eNaZdb0jEVEsdJwBnH2QMI
phoOsG+Mk11M3RhS7JIt8dbeCEXHaV0vNXToAsWPwLFguyoiYVXxXFe/XnRU+tMi
t6nSJXatDy+GQCB5227fLP7FNoSyfMmEPWUJ9RkFDk7/oAqk+jkGwg8T/O69a5P3
q8LI7OPlYsHGamQESe/KPToF3LH50TSytZ77UKjJthU3L6bwZiTNjcw/6WNgNuzg
3+SXrHE3IsLgaZOYIKu8rF0EFpLzMwIDram29hvdqL+goha2e2jFJnxHivv6vroT
yB9CZkIaIsR2ze/sJ9zTyXWRExys6wNyc00cCmCGRQ14lecDmyk6yGu6Yinjg2Ok
InyRMSJPDo9OPq7ExfR4hhiyNN0LOspWaMlu48TSBP4p6bj2Wtz8MJrLOzmTntNO
zFBTtKEk13maRxWPr6kO/Ga6hmzKfatT2agzSkOh65TCcAa+IQ5DlFMg5f8SF1YP
PUAmNtw2lSsm+CBvs9dKRjERwUTv3ZXHgJnKRsdHf4jdeYy6hswQVyFWCYYYJRnq
o5ou/fL6a6oIwdGOKUFVmKC+KPLd/Cil7bZVr0t9VaYrpgjfBGxFIhviLLypXB1l
HujqB0cEYBC8DjxvaSGxe74aOTAxnJKl4rQIEbxUfNaaXqfi5YNZdgS6a/LFRwf1
Hp+rpuWQrxZji9mQ73PedDHA7++LycxWbHNutfygDjlLuVPWKYwU7C67pL6oscNo
0UnNS9q1ya6cQNtYy7rMTu9LhZVTmmhCCbJ4MuVAFBgzVPSwYxhA+rWNyFMCv05i
ppLIZblceujFyFfl2vn1f1NOiZijsgRs57YaBEPQWPDGtMXF8i1ZNMY7cGvsQ0af
QAyLUFPU5aKK8cC8k9hGLQFvvZuTM8/Qiluq/VzPuFArSWj9x9q/Wv1Mf5xqyR3x
eO+MbvQah7IvosXyAMJRwNfXg/P2csT0XXjc/sXN/i+MnREYN7o+O/tsK3qVI47k
PcJ+swdJSfA3WL3OqvI03L95jGjjJJWuarCYc91KXu11kiRicvXma+0pEAez71do
mCO74WIFGKWObfYEc5J5bR3hAO2qG2VIYT2KuT8HZuc51yTyps0wjV/1worzBG4G
+7ZpSv/ECjLjZsVaBI3Kh42WPScF8YoKWEcvbWx4N++If3sOww9qPLQCICWwtdIg
vh5lk3D8J+fZOMDE410s0yXC8fUv1syJxCzUAbi9zcNnaVz1jm4Fg9MmzeAZ/Oos
jiYoBLIh+waya7W315g7xxM/XKnnI6DjjIdzvbjx5/gpkt8+mMgzamlPzBAoWGf4
0+eEHqoVtktpPC9cWGSBulrg7O8JIuoZGW4oyea1DiqJU7HbyHmYiKkQ6yg6XFeN
IOHOOUdLUlm/Es80sXun3AdxjbyRYBbIzC6n8Mlx9QE6geBvnh72ds2Rt8BruHJc
luEpsU+P9cO/gA42gKF6TzqZbz5UlFNw8p3QyKsEMRsjltbzmt2BDnRqbkZIa896
AZUt5J77fpP+mgTrcwC08ChTeU4eZEJ5/QVsw1tmN/gFscw90Kevjn1kUGYUKGCd
x+o41q7dXJq09ECugcuRrfPzNbfJGrNjvWrFr6KXjFLr2gOhPQuiOzG1s3gjKnfr
Dz1hZiGLUuIYXJT90R3ZJmOIaoTSl+qOfLk1o85oIYhCefm/TNUU6sB8JQ+aGQAw
OaGzmsY1Uy7BpfaT3bvZKl6Ri1wZt2w1Vd9Oe1C+1E6D3iRPKT3r0K1zaL1sPojx
RvCdcLjt5YchDyW8qH0cV4njDj7AESmQ7SSzhFZId7K0g7XhxovC/Q1lCby+OYTP
u1S0TK8FJpRwIC3h9Dwd3xrA1/XigtXK9UFA0rlyCpp06xGLWmVqhbODdxDhzm+M
t65lO/1wz5vLP0e6ROXIwR1LIKoccxJBTPXUtgHox9ItwpbR3VJGbVtE35c5zzqn
MVPzkcseBNsxbgruwftMFsj41vyGJ6RAA2yrLy+28YvXzBScju17Qda8A/+4lWAX
AG1TNo8CA/kJ8uQRXh7Dr5q5g2wloVhCdH5KSfpBUpv0TOMnjOTleokiVEhlXnld
kxJo3rCKGNjzIVibI/zEv/J9jP6rkZ/2YP3WJ8nowVu2FKecHFV+PdGbNq2X0SJG
Da4taFehTKY6twy0dg1ffgwjAo+9OnBYpUuXOAPqGkMM+MQeswFICGQGDFPukF2r
SN+9YNmakL+gvKrzm6E5pUgjjJe1+Yot4Pvl873gzz1xqaRf6Ca/4LxDqmPy3HuR
u7tfEg/n+DynA9+rl6OLxSvSQO3WJoJteAEpTRDoMDPzHKzmu/vFwHye0qRcs6Yg
+G3E3E9NNIXcbusRjWM1CJUAONMUSus9U9Onx7yVeYEQFAiIVWBQzwvqHAxZy/+G
PFxtCjNZiwazkGkE0cu/cs9Hdot2BmWWEXU1NV1knQdXEFNX6vZA/KBkE1pRcj0D
u4mLutWBsWki2E0AUakUsx0x+I7dIUtOSzUA2aThs3rIsWS7Jj+CzvnHqs+jLgSO
mCWpxcVGo3AhLdLSzDQ20//O6r2NYDhFBOE/QuJSd4x1oRvPtXqBCmMPBtnyuWJG
YONoxik36PQX9auqRUc88ERW6NPlNdPHVhNRuSLaJPaDQgB8tQMH3+XUAMAOgmsK
qxp+yBOqZRIw5u5K8KnG8sl1asLWVTnDTugdL/Acs3ysU7TkCypQo6OLu2YfVtJF
GrX3XVFa33+DBH6i9R4u79HkBT/NYcGCK4+9C32i8+hlnmfToztRTN8bY10FM8ij
AQc7L68p7ZIfMWmHrQJn7+Y9N42dMO+yjHMdBHRKsdJXAoL6KiiXAZrIOSKYuKHF
AjcOyj+QDaQfn/qWGokQVgDG9tcJ0ceNYWzzDnEHxznaAjLDCCPIzYeSFNxbcO+w
HGeoEGrJKa/gDH4/4h+Cmz9LXrP3SwCCfxDXS/tuzrw2MbFXh48arUdp047Fpnhb
Kfpx0Ouz9+suiFipZjT9dB/9fHCLnHg7SyVcsXtp3HtaY/Hgvqi0mZPrAySzFQhY
gdvwAOsVlkpmBB7rGCAsOlRMtp7TsKtayDs3Jm63Rx6f7LTON/5MMKcbH5nPOgJv
2OwGfvsisbDxh+c4msnkV4nNTZiKZ7mOVPNu1X6ry0IiKAjd30X8X17fQuPj4nIq
I7hWaeI1rtdoOcPyYDZcAEXS0F6G9qO+eXD5lho5Mjk8mbPl7vztneE/YPbvV4dc
8t87IOUor25dYyXQ6hNBQPM87y6laYq02c8XW+aEGircujPLJ0j2xcK0vfuFL4x6
+kKb+W0vnsgnD/P50UWG7VwNsrAK3WSJzU0jmqIh4lpOxNhugmwreciEWiujpfOK
uvSBZbWZmrgQo/fyjlqmDH40+LUDkxaC2bZq0Zg1ftmCnkOy86bNq3H+Jq1xQiTQ
q9paNku8vkT6SJEdGwDMuSZAZ+MJLaONwQ4rcUANMdMapW7j9DdcwN/EMep0sk4b
sCFWbvaUcMvtM2KQMWaPge078RI97AM0Hf9dQCUjGxVaZaWVzSRr4QuYRQ9MLakJ
Mnvk48DLXqzlfFGspFepySrdKOmH2U2QAYSfW7YFo91t6t5fAh2sx2+gWHvwwFc0
/wTOQnRx/j0iOGVI9DRsKstpT5UpQBng3xTQbKDF2jUjR7yFBjDVpD+O2ZawH3EN
3tP4ZnV0G05UjIJF4dTo/kJz8HhX92/luwgrCYfCw/RK0zB2i0W3Kih8L87pP9dc
KxgVGmDvjpHxGh30utDfTmWxzdDC8mQzORZqfnI/Y5syge/8UYnHVfv6jC1g4Kov
Udfeu+uK89gsFkQgfXqATKv+amX0z3fu7/gGdrrtcVAUXD/ZOgmyryZHbASxt5SL
u2V0jxhwzT1n3hmvyN4I8mUlOe8odlVz2LoQ6ujr4ahDMnVDPL5GXLQRdmGZ1skj
26VmEQ7hueCsm34lsu3g/2cpXE/oZxYEuXzIelsD/eoTSBwKa8sE3wIsZtiLxaDh
W2ioCg6Spzl/KUu+hm/n7tkthvUmm/naWNwX7nZ8AEIk/qO9j+J/P7I7YT2+SjCi
cpmLFA/dAtn1G40Y9lb/6mwBXjV3XaXUPwUK5EfwNPffIriNl0HlFUNa1AFZyPtF
GcVVIVm2w++BT14Qmpix3y4m4bkBfbhr8v88J5AtYVySsJQEeNj9EwhvjPEwXxOM
h3Vqha5VOPfBwLYlsISlweHlwZoBA4abgPcFMKkwBKcVvSnvgUfvBcw3OHewxORK
w7z3rChgmS7l/A25pr1PRbsjaTR/3988I7UbnNyRK6vVgVmSMF1hqkIPKcYXTdkb
Z50ARn4vT7ApPaKMPJ22G5YUg0BvGQyLQjTU49lLUOL87/Z4qcfIYIjdLd9gxzVU
TOQ6IihlmeU0K/pzCUSny3vCNyYhc6LcE5C9TaWrgjIbKWNOpAo1zZrJkidC/vBq
gwcLaxlb1kvnlS2U1UmXT6XwZar50XPf+wJM4J+Zm2Sp5OCvQSv+z22o+Vq4aJkp
tLEKrnBdmLUtnKZS00d/KQH5WVDgymqG74XGN0P/v9O8qzfu/+17daTEaQgwuBuJ
DKFOKSq+7wmYjhOGiP97AASwbp4GLKrQTP51pIhm3TM8QPQ+wlAxfhdGyY8lXZyE
hn3BwXvOMFjG9N95swxuekOmC5c8IHYTEqa4hybRTub3HnPjvHXa1aPwS02O3ZG7
re+wc0FekSC6C4wwNFgqGF3eyzvKCWw8Bl47Ce+XDYWjTlF5rCFJSsD2N18xoHbH
3DW3Ohppn8BridqlDUlnQoCnWvOci168zJFCpV0RuchU9z95OZsnDQFmp4t2BqR+
bWcsDU0ID+AYLj74G8k8o5vmKvssO+DuGH/8XVSqxEd4kMRzgB7aHsKh4ZC+d6XL
GoFcx/pWnRoyPnnC31w038DL7IooD8J7hZhcZyGIpKV0Us+aE8aFosOZ4vVF5dx6
f4IvQN/KPcRzY2pG7lGFo3HeUBdXZe30UC3ktQG1X0NUhB2sXnCpkf6+n3Y+JzN5
QqUXQ9uZrvGCVeT932gfM2/K1iX+g/wz8L6wILs7lRSF+nFy35rM8mb0Zm/wOSxH
30etZ2od3DRCRliZdmzSu9vb6DyYP3M9xZnbbWIMt/crmE4NGF3CZurW7BbTDkVp
OG/yUw+GM5ikDdMwG1qH0knCPEStaHyVzx6GcUn3r9Nf3xBr95gjoluDsAEevpyy
XfjQ2CmwM7UvJfz/sDSQBh0Cp9z9tncsgsuq371dceHn1h931Xo+ed/4x1UagWxR
Glg9tEUAWAbmBp9u6F1/X8DeNO5jgzWO7TI2TFSsZEMJ5djep1kXOaAwLhu0owyX
4GdxT4Nwy1orFwFx+rhgTcgN6II8CMCiyEmlaq+nJwk7Ih2+aUWrhiMkcrQ66waR
4hSfpxY256/fObgZYIhyRu5ZS1RSwt0T6+sh0HsQTzUsM4SfvTL6d871C5n+qEFo
rZQF3Ax41baG8A0Q7kR5AeUuMOzPaEMYAUGPuOxUcpAgTv4ASzM5WNVpDbxRtp00
q5m5gZf39dowbGG91m9IeQpTaoJ0VAltKTJD8iiu3xE2VSjmZq6JDWdw8cGJpLIe
WZ+mlwOyUq/T6ufBHs1a8tzYfoxJyKN/poeaaetyeyjI91Ika+Eu4Lv9XVB0S2jj
SFuLbMoXDuiGTxx1TFF7NGW1rBYwJgnVEvom2U1tuREf4I6LZ48YQyEtS9yzal6L
fXWqvZ1+mfzQrNKo62ksiFHM4HhXDy86r5V8zPiy7S73DtRlaoq4N+ULZN3vEsHP
TqwrOLQDddQcJnf8ZfsZ8Stp8336pZei0nLFfqqFr00l2OOHWkKZkc96WJVvwLXb
zz5gKjB8PvHlsd3nasJ0X46tP9UQw6IouvhqoNtKz9GP8Y3lpCW8GUmbzO09LX/y
zlzkdA5vHamQ+sGL5oypZ4dtqLr7Wv4wCBwWiYpccQuNfAkxkR2l9hjb41/wuQd/
9VJ0nz1KHC3SjRjETYtv2Esl3To5Z1GUYHDnv97dnKLOJiLcXA/GlNnOg6uPNqGa
Ic4N7JtL77VUtpmCgpzTAubXDNsmDE5bhD4tN4Lqtxud1W2QKIxNXUvchhzdVqm4
Gp5y0EYpjxJm1MO+ZJBX4SjEqgFQgBYGH1N17epeOmC8FPGxlULvf6N2TZPTsMG3
3KoO1gbWa6wFvJDt3CEgvY8sAc0XjoJ1NVHaXNNlp6afKtVL4baUCIyvi236kJXl
VkXpGqFrXblAFen0iIg5qqfS06e78ugZH9qKKyVlcVifgdOKm0A5goBrDIZZNTxg
wL40mn9Vpa1FBnXUMoEkp6Cx8ICKHGCTHJ7OXF12dd/Eu0ztihodGWFFCvyUiGSQ
BUTqvVp8+vKUT/eGG45l6qA3e1y45LqS0B0x+ZofwUh1vswbDrvWWWbZ31i488Ja
/4vFOwrTA/UrUf3gKT5YgsBvxHkbTWOoW8a/xPaa91hfFq28hjaxCQMRDiVwX9zV
6ot6aa3QeiU7RZ7sQHtWVjYCOk/zMxC6sACoC4JD+2nq7i7QcO20GFwnsoBevn0z
g6zy/MqPdHjMOoIIf6LjoFpZoIUSi/9qtOLnFEIhrL35WpHi+17WLWCvfZtB7f74
66mjPcV7UXTfmESJX+aFntYmcRm8m1OH26/eLlKsX3LYruiovOe/RZY6Yd76E3RN
0U04eqrjopMmPxVv3zH1zzcUFN5wYyYSqgVYzp/u5IfXlGNCixlza6a+y/GbevxQ
jMPujtie+/qGhW7o2hFu4miqBIi1jDbMqVOatQpjZzhEOJ0MWTMV72RXe/VTBByE
7jCNtjsTWt3lK6aIwGoBJjkGAy55vOjvQs7cwd76A21CCIbW5I543U0P/I31zhZu
knKE/+d8ugzZbSmjpgwqywV9/RHuP/mr8IHef5lZMtwP1e/wkruN35GzjN/vsrid
ByszYmALVFdTYMIych6TpAD9EKFFjVIcDv2tUg0ZtkKJa6js4BBOYPNkvzjV1bOI
u15bSPyEvI3Wkt25PrkGjsiy9Kd3niosKuB/zfyHyqukIpFGDWFNacilw7ev7AlM
ta0FWKqykw9YNKnFxhfyaHlap0zMkxlKdkLJ31wXtXotGICLE+HXJc8sBqI0U0mu
DL0wVVX/fh7F2eYez4NsmBdcJUHplGmqy/NSYGkcrGZKwRzx819XtZgkbC2aFP4S
5L0gE02U4yUMXWYJFef6jrSBTwyU7XL13L5HrXcfTiWfluk4IC/tDp19bsjoiPQU
q+LUDnMsEe615+S+ZPAf4hw/joNz1MJSqjD278q5HirrGvYJ0KN8thfAo+GFhfdP
P/rc4bAiDDCX5prSxoc8LcB7l71+BAR8Dc8klbFOmuJ92UGsOwcDqNedqvOjnuIK
LnkVG42YzBEOziqdA2rg6nNJhsfUlWFl4QEDUZzpVsn9ixjimotBMqqlLfjOiW34
no590onVoIIA7SCXuZ+urQDznVNGDFyOV3XrPHXYTVJgwUQXDLhxTbAlnQEZ9W3V
Mi9D8tLu8//R3fyVrGdwO/wiNFohxYUryPSdMAMYbgI69U17mJ1UQY8HTbfq0l71
NXH8nd093cq950dGm7PUF6W7OyBDbhzFaVrPqqeXG9U0aVcsOMoPhASMbPUkUPM8
RbWzlxbvpXziTlokdnLRcgJ3wKpR61KqHVZU1g4WlyVTEayJbS8vWAVchjeapsGK
+SU6yxebO7GBlIr/XpRiwBdV+4nt4iLqzXdxCvXPRRIplv0y0+RlXpvoHfMgVy9n
k57ZpKIgo+jPZJcbtFcBalbTEIaR6buwWcdwnNJ9woZiN+K8k4v47Y283p9ah56k
9TgOahdKVejvhLLvQSsBX0nR9NvDFHk4hwEeWAUP1zk62QbRiwEXBj9HOfkscQtK
3BNFWyfR8sFN+MXyRYU18iWpdW7dAEeyEuGZwCGmnTlYTvd4jw/Bwnj5wcBSM6x9
LW9tF+TT5XgJ2cdPYjqXGqPjySYzjM6/JumIPfz0ctwP4q0WepzT/oTgtxTFF65i
kRk5EB7myqkjH9KuLpv479RB8ajMPoL8tVcld5BcXaS5gyUR/MJglAbeDO9ZE5ie
oe7Ee0pk1EV4ltOoFHVc/P2L8qSItpSOUj9vAmivqBhGVVx0oldBMGFbQevVQz2u
gPcA3AK6accoOxuYDx6uMW7lWUgNxcAOabYm9n7ykH3a6kdD9INsm5lzQrMwVWks
10okZAT6bOVpXqpKo1kaq+iKtk+dYuUSnyIL3OgEtaJQt7H3JIjs4kjzHY1DtgXh
yGL8Uy1J2mn4x7cqtdmCoOutYXWOxD6lYJ3KC+vM7LjbgBnmZuaoPVAFIzmb+fgu
BS4BPQVj/jYlDTkoWv/wiCAilOXEwq0BLhp/s3AIUVP7vqTXLlGcnon1ZFa5eABz
yZK1oP1ihEwLi8A0pFzWjt5thCXFqb4AJIS41BFASOtVhKXUFNMbx5f99Q8xOPVd
/gfynZIkGk64bHUMnVjXlRpaNCGM23+rXnRpDu5755xCkSFzA2mxoXebYv9Bkqw1
RZbVeXsqq/sJKIYiDCL/H1LrEf0cy/7b/MXqAA7c7CpbddQGuOdxT2Ok1IInE1wL
l43ZeqCS51R6wk6BX0AAviJDOKVlgvCNn/Xs05jLVf1r6cZHGNCuYd2q/OFEr7/N
pHdSr0DZRFwFBhfUoritZRTlukFVwwJVMTkZ8LcjkeemSDSgo74iC3IHxaSweugJ
DWNyQZSv8pzIymxJKhARpiHSyTrYpACTILCRHPPF7zLwVkxsOS4pk53uBhyEU89K
hhFWkwdILIkoSYHRYDhkv786gN5amPJ3a+pbT6G05dZTVmtUXL+OHWfNpyR/mVO+
/Q/bQ1btAXX/NcpqYx1raN+tN4f8VoswFsCGHWq1r3T5PIRLFX12KaL/OxLvPhvk
QWe2GV7HZtzQl1dHAfJ7XzT9y5j9c/cQjtqgySXNInjUE1sRV6mga6BYV444Tzmv
8mUbSLmvyBNRkuUnLXPt/o5OuD8j4A15TTBZhyjU5pxF1IVWabbrwEF7Z1VP54LR
eESF1v/yLb+InjhTjcmEBMzGeq90wnU2e4F83cYlcr7uqD+/ZTQ9v+NcQnNGUKwR
TdTKUpxyg7RWQQMMUWpRrNjq+lkbu66XwoEOPB49Qfprak99hFZI6481s9ZXy1YP
YGLBYEkgVdWYbbQkwud4FuO8QZiLEongAJX9M7K7Dw4b6lggThRFIETJQmdCkkkd
lvYcoH86CYO7RQzWqwBDF3DpOdkZxyriNDvQWZST3BGcKuuMnOjhQyP1inK5XXD+
BUB59pBA2HRRI8GFTo6TFq8e9GFRFGGV1SzPz37kxShdXqQ2hoc87HvExC7Kwdzo
ofCu7tZ0TWjGqdeVyAoDbH1sxAdgWe24jMP98qwN5OA5JHMsF6d9gFjch1gsUJ2l
50Ybk/cbroD92xyz5wtO2rCWBXnHodlRuD7dSEmmpyg5XIinHqdvlE1lKX+bLVHL
HjPQOVkItR26TURG1DjWGKbzrdhuaDLN1CjwlkN5t9oca+awO4W3UTtUdTxKH1/1
TO5sPms4+/7Ht79Jhi5F8vvbWajwmIhNASWv6IRdvIESQE/CIfnAyKtZXce1Daxm
RGpAEoS6WV6u9eCXkSSH4/fOKs8sSDwK9RNdDlTQmWPC2jGczZbrgeVbBpwMjJLJ
uHI9XXr273f9pfQXOhFwt1AIHYxJdoU5Zl+bVKrHkqpcxO+lEvJQC5z64OLYV3mo
lSgHPElfOAzJVk2tYPka/3Y4Kzd3v/+RT1cBPPrvctvxxq8FTA5nujweTAzGuAsr
bi+s9dW5EfFR8zqm2i+gGjI9HHJQB1ofzbUoV3OFgLSfR6MI7+0wgtZNcggXjTd2
yHdZLvoCm0YrSh9RqQNSNCEJ9+vTZKMKoWkX1hY+MZ0yffKz0vul4yVRowfISL2F
XsY+d0jv4iMZfWhdI/b7jBdcSg4qpCospRWFMfxJnKAvIniL3pMzW3iCR1ztIkoQ
FcNmrS2dml7myWhFLbCKZOm5OBmybwSVXOMUHu3GQ5ebt2M7Lcj2j/YAngG6oTab
+OCV4Or/WdSId9L/6nno2y+kuse+vIyrrCuQAz+lKtXitNncAklnzAbqppeYomlR
Hgxhg4h5DhnDM5jXRGZLvU3gcACl4/r+xl6VxqTRlC3d1Dz1t68xDKjOq+A6ZpI7
g4douzGhowX0lfcddg4i4QBriQ7cB/Z8l/M/ti7Qin9Hn+7w5G1sVN8ogL0e/ZDx
nEK818XQEhmskoQ+pr1fe+Uh5R7KiymUBmtGz11mTS0pjDX2yjt+y7hKNfK30sir
Y6XHomC91luVaU8QeBmRRAb7Gq1xbxBlqHUmU+IkRTAzb5gNJMHab3jca0apkpia
MODVKPeFrWWe19ecWXkwIZo8fCuYHXsMWwneVqbaBPoCa8QPHMqEKfqO5+XgGPso
YyPDmpel7UiOcoL2AnmW2OSx2Hi/Zt0uX6Ca28SbpHbUIVTie0/SrSA70wWZV0IC
kU0GrKwRCu7Hoig/ql04xUBCrT4uOh4JyH2AVDDCWTbkepX+RZavnGFIarbyGG/F
wHrR5iIULAauIJ17IbXVS+2/cQ9QfAF63UioD7M+WnqwMLNQwTd2x4O4g7YMThnY
ooCpp+x83ubrJqNIMcQSTibDNZtaipEplEbrFYruUCrbr7VGBKVO62VP5p60olxD
WEupZ8p9JZHAXWYhvt1ZNYFgMTcy7dBo++/H/dccsq4Vborg8Fd5BRoeyV7St7LA
AUDNC0Es6Eq2Wp+uX2qe7Y6cr/AMpAv3GXtxmvGmEmWm0QM1W9I5mXNXMJFmrnrc
E5uwIQt4s/fSfarxQU4BIRos63Og2oICU/Qz6KZSWBQcCZ/tJQvf/s6jMmAnPQ3Z
qNorc4MgcbWMjbbqr8fv5Dd53VF9hfoDBzsGQ7Q/NiAdwARv70HyWCReIZHarZrC
aUdsrB6X9lXwQ3WG5nlUaCC9bMbmcG0a+BGYnrSOnF73IIM4Sl8mzbYWdST0HUjt
mcJHTfrAamJy8j6t2oEpuMfJE5tPKfkWesb1G7x2NoHj1qXaDU/mhIACo8fvOcRY
k8gm8YPZLces7CYtMiluGxJJvTnvTc5Fc16vhN8/kuW3Z7au9mWN8DToVCJJEDV7
PMQl508mIdWlkp/FnaXQLtoizZJKG6wWD70WHEYdU+rCIf0FwvvcrCEgc2/cHK9N
M0kC9tKrSxSG8rAnPE0UvWCkQ7f13UFfE4UjQe5c498EOM1GibTMLZ1+PbnHbAPb
mFJqK54VC/lxmaTY6HxHmtPaqraQHshxYPE506h9FrKKRLmkvZKKOgb8P2Mg8u7v
nVVcMPRg5c0h/EivPfGX5KMVYrhYsVXgC0a1pVh/gGoDDgI+1+gI7KaDsX0B1b9y
MonyOrPOwDeN4bU20xnmX0/WwnXYjVnMm8dB2/aX9uIxB1A78kN5fRcd64ActZES
/OGJLLNcQQxMdfVKO4AKO0R2W3aCgcrN0FBAPicQuSBYt6WITXc3vZzK5AONwLzT
kAJly7NE8fS7pe/CJU+xMWr8+OCeVcxt/ZsRtDT/hwmsRT7ffGc5AGdEBYDZ0EU7
TnrkZ5IwLP3eUI1Fe6Pdv9iIC5Mc2sLKShprI3bqPdHuXvbKE53XM+nCYHdeAX7/
iqh43bWX4lOj7ObGGm5aKXILcyd28KlYW+Uosa9DgbAQEWSx657T/VlZiifRpQOq
FdO6E10CtHhofP/+mbb7ksvUgWG4yKbDMdheYTUEowxBQ3EI1ryFjdef74UVzwCE
A4E/CeTr5HXONYWz8fyueZcshVb1TxZJ+oqrjnda0/zHseerDl1sugpa7FDxrZSf
IMtG9n5RbxbY8JO8KKawdvT/EeMHkzmpTYex4N76IR3gMFMTC9JSIA6mtVCchFgX
E6K0HJuPW4cGQD94xQI5rMP6GLxcFV+mGN5gI7jiVgbj8OCaHJ75bKKArzDa6A4J
gzUeSj+Vx2dtmdY7sa2KZ8IEY0EmeIJTo5opWzZ+kHyqnPOktPBh3g9zRBuljf/r
JWIeaVfuvSI8hGXhoyUf1dPxwjxdiy0HrenRBnGQMg8A60D6wekq8pKpVKuDBzvu
bAlyUglS4qs5f4/rzHdF1m3oAhR5UVovxyOPqAnWqIUqlDl7GlwBaJGWGmTeANSO
1o6B4A7Rj3NHwFMLndeUb9ZOQpFRx963ffAGiWbWlie+X5cVq4YgiB38IO/JtaqC
4PACfq3mHRLYSJ0llXZulCei+W83HmtNVYPiU4ivUOxj5Nd96rd7qJPCNdih65xq
gIxf34bgcZxKfxVUDm7V0wnxzY1l4g4b5Ae/2p6YXGglT2+nAojvUZFmFYiJQ8WH
lJmXbPsVY+au5PuVSoIdvM3I62qNrGZM62gC9v0Ht63iHlGC5dwdLwcLXhAZChO2
3YiZrgmr2bM+Aro5ZoRcqjRaMhWlX5dGca+Iu7psMKr+0eGKqEzX9OyC5kLjQ0zb
QCoKqSfeaqlATabYOnf7eSgKfor1ZcC4SZOq8tGbAWa2nNZKY1Dwa92jIGAFsCr+
V/VV+SE/qcJeDvWGAghY9oPd5eF33HCmtLjExcOZN4jkkwPMCf8LWLJvCvh4MecO
cbrVNwb4/wOjju5CKfKKNEDRokDJ+aIOVTRXvGMlHT+V+UHpyz7pQZ2t1xMEFbX5
gwrWxif5CxhKF/LgvxPchLcDbPsZXXBhWFkF9nY5oDaTNbg8KdJ6MjvWQETYGgBs
h+BvtznBRYAXtFUjS2fUFmvDWVmS4mxJBE4inuR5MGfrM0CbzcxoSEk5gKZPhVmk
NVo+JffBvUcuxDqJxpoSg5XTk5UiDquOl3+D2hjDvSvg4qd9Ty70ZY9UGkELJySs
Gc60hC63mKxlDYYqN+69dsrVT2Pgv+NEkenPu0eEObzdl8qLlcaN0NYmwdfr1NB/
KbrJV18lf9v2ARXikgrsFiFVR1Tb1FPB8OXjGjzShBYkJu+T3gTil9WsNVgE9QYO
bkScBVIpYMkHdzv2Iz25W0XKIopzWWouC3s7k1BGqjsTG+7njxMJGHJVKLhUX/eX
exzNQaT2c7R62Bx4O/sW82EiMuCZVTn6I6pOYequsrUNpDcgtYRSuHu0P70YLoRV
oPiQoL7Hcs7DK0UEH4a4FzO4ipc9g374mJWAvrggQaJaQ4yPA6NvhgvJLB2AWeH6
rNkssxnXxJRpI8jfw5CXZBkqmpgyX66fE6O89oT+2nTdTDwSPLpDcRVfDDekBr9T
v3joi2/6ly8/SbmeyhJC8SFIkEhtt5uDjHaWInn53KoqNMz1gEYWEKGP35aoL1rp
zMRbKUApp6rT3CHqXIyCmwxYcLJRhaYNqWkfiKCXMe1gQjmRO95RCTUH6gjQumsn
3MiSu3nWWeVkq3PN1REGnW7/w04Q4kC7JwlkY8mLMKMpje0IeBYEL6o3H7ABv07L
r5eP3H+zgnEEoQKc9AeY/6g2fqrgaFDjo3yph+MzRhGkXHG1emDMba94cQY1CK3z
oiUtm5pg7EHLfv9e0V01Eq5sT9LJTmgbOnvhhlRkNNPErsjkBC5SbBsCBcXxF+H+
rzwGqhLpwpVdqD4Qdt1lFeqrQauPCTWqW6eeaFFgGXEurzjAE0WIJWYEGQEeQDSU
8PGLtoolISIneca8XlzujMtrr2p+wFYkxPqmus1SzLS8JxP81q3Asw9+FVuLhWSH
CENazpLEmvIFgcyBD1RST5m57wYQb9arTmdbHOtz8Kvlkuj8xKRZzrzKUbiUZXxq
JwI+88LswLtdwNPLiog0DRFZvN1LMX5oKJNrV8sI+a+SD8Ju6zaJKCbaqqy4kwqx
MNRkC4P1/ATOKeXyHLKkpDOLhv/Pkhlys7Y+WJmZpmsG9+sd8IAiTD0ri2VA34hI
rR5GQ/ZjkGISf1aEuBzB/BFLCTkpzqKDb1+LTojTeamTqNNVpkAWVxvwjwWVvYdl
czv9g6pLR79br25o0o/0y4w198sukwevsuycrNwZ+A7ud848+tDbHIhZmu9MixIg
6gPycQ2qVlEaOBBiSnCqtFJqoiA53UafmGkZg7+tWNXBGqGEJWlM70+pPtl+IQBr
UxXphXkfZYAZhbexcRRD6vN4zuOz/AC4YY3Ki+1zg48a5ochCyNDROzE/wIhLg68
KGAUl4QTU6JZoSh5nesC+Jfr/tSM9RpaucUfVFsbikqkx5d+WxABRkPK/wvsZuSo
0x2d2pamVysMSpL/ZC/+G7kuM5E96f3G5AK+rw5r4Om0h18dyn5IXoGBz//6O9fd
EzijT0AbqquBZNmfaN3VGNtfsRCxp7YWq0HEiNApiJYXGQgI45W2FfqE2guFS+9G
kirZtEZE5k4Bim/Lqg3LlCY0VsBDD1HynjojIIIkayU3xYPYsUlPggyRfo//9i1Q
xvhkLsOPvMu72ALJTc/irJKBsRRW3H4nMoeK0LVODBySAI10qNxRS32T3m+HChpC
dy9hTKmdD/JAV4mnVzxaqrjJVRobhyxa+GDDfSqUnrI1z98wl0uhpkJVEUyuwuLS
1456CijShtQN8LZfsY5bLBA/AEJ4uFKcIxd8bHgCYmeQvsbo7/20ZnLnIxAXEQfH
9psFwv1dWAChEopK9KwpmFeeEfEGLKvTZ8aqBXlLmyBCQ880/48TZ7dlYbtvzAFR
AqarfryLaFqHLHV5PKuQKB/xNaOezyBW6rhYJgrRvpkLcM3pfLUwQLm0v4YsYXlN
W0KKnojhfdbRVGqX7Bdcp70lvHMVYWOaNnl8qe+1sQdh6fw3RI9M5Mx7tRq7XiKx
V2MqvkBjIPHNz3UWZC6Tq3JxFTfVN64nW3ipxvkjTH0VmYxAJXpwA/+Y0eX3GERt
Z2QBiYKZkYxNCEhhCFjOWmW6Jj1th9xuzLP2Mzc1oG+3lWpDPjJmorENCeHI91sY
VMdMjFFvo8Sn829ofzKglyKy9c5AYhjKgwBJ7tk2xDqxXlnOt25ZpIxpwug9DJnq
Z6ZwJ3fWcrLfEU/6EKH2Nst4FqiVX/GlHNUV7KIvOaxYNqKmK9g/l9/XBTTxChT5
yk1PA7652HkmC6bGidIgMYnxjh/F1zq9leH5dNKHq8NzPD4QTngsS4D86Miejv2m
z7Q1FsB7SvO3Y86ygaCAwfVFwi3t8hXbqjIYD9WRYnl9Rxdm/WZv44HEftKb5prc
Yb2PHaXyVcjsbsFcSTrB5XbiqrNh8dtHQuqLi2/V2wxwwvnEu5+fWwTN7TSqmtRI
bakqLui5aD7w1/O8FgwjDd8gxw+Ua40BKnRGyakuO9BZ9HB8TodvWQLP+hqtH/6j
8us/HAahZpy+DreBdqd3mod3ktuN9LeK/S4vYUYGSBqTD7gEIVUbdkOZIRoKphEP
PmaGwbb6yZ5QWI2yxujtSLTKG72+ETjEevV5+91WaAmgNQ2gx/JNhHkt37yEfIS4
QFflzqET5wntTigZOudMXfis1Z0JlS2rvoN586ELzDfk4LjypVbtQQHgn/5U5YWr
Fi5M97V4iHA5p9t2poxvS2r9hKSW5tlF0gQTEPWXzcmXthSZqVU4nNJ4Qa/zK61v
CRwIISeTWbSH7XLQjeJBf4fh25DEokr2HU8cKWk6wD1VzYEs7zBz6RzXfbb0pb9x
lsNQ1SA+qJA39feAqn6THglt7H2eK28FLAuSeFB4RKd90/eM8g5dk+nlVYS7U4Ih
ZRXYKEMlzGTczTfhKX7wg/8Na8UdEqBE9HOXOJnMYquSgx6h5w7Iro8x8ws2zL/1
16uy/j2IQ2pxd5S7q1XpdW6n1KeI9Oby9irN0lDOrDDaoIkMCS1bqcM2t4mcm1vt
9GMLneX3KO0KZT7HQ/mN4TQc4z1DYUIkBspxzd/joZ+pP5txpbnO/kxJrIyXiEyj
DFbUHRZ7f+hdmWkNEMU013yhyfeg2D/S6beMo3uSMf+0YOBnTPhORVO3TKPUmWhq
rqBxnUDPMJP+kkXWGrGfJdrCgl9tZVYSIrfPg+71SUWNYjc/a9O9wV6EocrcNWNZ
qIa9maQjWCfVsz+iDnU0TL7+9bV84E9PHtMiqzzhyCbb18cni7of/giXCBUyIfwH
aOLm1etOH4ljxXFEJX6oQA7zFg49heWE7VOLNHGmnFLcI/zWfQzyc31ga8OvGBi7
n9foGxOx1GvOsWOw0qNT4pNRh2BwcM0J1ejAtXp6xzyGlrPhH/xttt15z9zpvnM7
p0be0pUElSNCbLhy6FXXbceIgBwalrcoBM3lx2jjyVFvKL/Pf3jK5Eu3KeYQ2XTN
DJ/JYINt+zPCBAec3mRzQH90x007MD74Zat7IBRLi8x2h/dFCxdhbjaxddHQu6Nk
o4cM1sHQM7Ct6f9hEoXbIn/QRtgEbUGu3NuMYrYaTKzTvXyPsjDhlKJ2cXa6r/TY
P5uJ8vYrklb2Dhc/cylQRpGL9pvC9jcVGMRiZGgtb+Ec8FojH1kcbTBHddCsQoHw
t9LQbaXCHizw9VSnSINAXKjiVRspcnZlAEpx9flwzVtXQtJnRoj+jxUFKdbf7V7U
COr0OGc9NQEQGRfUMAlamgIBbwRQAPG/7NJ192kp/mHvETraEnxeyPVPlZopApVC
XUdhlU+7Hvz6yRl42tgrDhuA5TpkKvYlln+BCygvgSYOZ0QxuSEUEnXQpcGsJiE+
7/N8ehX18s1MGCfbmwPh36u7mssQrLqCyMuDQgpJNR5adn+by3KJo3ZtEnLHBeEL
w9lx2Jl6rqiG3wJSkI2WHGQcEPGEotoTCNWnpJQ9B1vMI+C/Y1usMypN0mJMG4jr
nu9rdeRN5uLalzpemrRo2SdVPSj0a1fr3eH8dBLf0M298l9Va7upre+cR4b8dq0k
Ovlo+Rmcl/rcOwFC/Gg3WmAomkyxvz/aJyHC5cVlI4F2Qom0VK1GvO+WvbBfgR4a
qZT0NOl0QbapWRnn0WcOq8Sk9mPqxnuTrTu2kOIpvHouBzKo8EDCV/Z9yDFMPuWp
GY6UzbFlZFEMzQDebmU9URFpbDiJHdw5usuoEKO9UJkyFrSANwoTzYDl62rhkc2i
tH0RX/e86CD9NP7ZP0rkk6PkwfMXpJ6MPgVDp3RoXvF/Y+sOgHl2eV/BvsvBG191
9DFtIwzG/V7TZkXSo5rqlhNVRWIQH2sScOIov7DyN4XCCvTqHEn5VvRH7dNT3LHP
z+I5JwPL86W8P132Ms1cdF6MzpTX9fQa+bKqE02IvQN9dVwPXhJWWXFmGBW1inZY
271rmaB/EDir3jr1+Yztx6oQUWEuw5OkfgvdlE4auj7QmyN/bkt8H/HgMFUlFoxt
aL6amtZJFtMBRIxXxfot3EgRD/aF9bjcqFh3LBJaays296l/jpfqWYmoF75HuSkp
2PDh8M7kl7N+bMfrIukhPMg/OA5xQcD+2dRAv2i9l7+GNtfF+ji2pYDrzEkEyeFh
EbLDAI0vX3Ce13fWdGW1Pbws8EvRS+QSOb68QxJP7uAOYEbiAnpXgsQlssAEL+dJ
91+vSURgXQLx3LaVEPFaOQIQa0Hygzx1/XaJOHAKTQn/EmFEuv+8nyglyXP47PJM
k0qe9XKVHcbHCtX5YBolIjdcHayTGuDF9UksLfTnbLYuq/6BPdEf2UV7BiJDjKKr
TtvwcU2tg1jP3M5WWDo/QfTpsL4r57xBaL4Gq1Cskewx+YLg8pu047ORj0eBxggU
Yzaclohp0x72SBg+JiOSL0nEt9NYL8ugKcWKX2X6t32DRlGdBvPs319RitGxo+DH
0MTCb5TXS4rP7tIV6bWtHilhZPLy6x0sWQpcmgi3KhzVp2oyd5Bsz3dtJLn8G7uN
UYeSBxzoq0wEfVqVS14DY0JEe09fIbu/pZGOEy0T5lmFhidOFaspd5EaWhpDook/
SQhUDoPUh3GtTOTQrMbmkrBgRLocHfng0iXYFzN7gkD1TLEJ92WFwq0xTwhijiiN
cU+qmH60XYxggBWmJTmaYdXYNRkPxQSLLjNVIYgP3U7niwFngdI4+TkvP+g1SqAJ
0Z6PVBAMwZm7h1tXgmLXDbIyET0tzQ4I5bnVcrh/iRFJIVVRttuap5BI3TWIMWzZ
uDEOR0wWjsnHswsphNpzVbRzivwo5Vysm/0dze0ZOXPUsHO9p4zvjGuHFDEYjY0g
vgOAwychL3HP6tBXWaCw1emmV5o6mFtbeinir+qXlR9SdnKcV/GPpCdZ49X+9FL3
IuRkm/0XEsTkR5U51B2QEOt/vXbB6/YtRwdrhZorMtsk0S6p1VnJfoZb/TWhxpcA
YzKsp8oq1VW/0PZ3BWzV8Cv7ajgaQQyGVqVq0Dav57rYPL38C6Lv4DtmGOOJl2Q7
RPB86nl32U+L6DaZLQrCGxCvlUywpttUdz+l3R35ccDTZsaxJDgB/1jHl9OriIcW
9E5B4KSyUBA02txAI22a4BFx6ETpRQrnztJy+2GeyzCkHq3hhL0YPOHw2VTbNQMu
KdjWXIG4dM5ZZphKafnRz/yYnZcBNXNxQItHvrmljf0hBwz8zNyr0jN/sA3ggSS1
bGVJd5GhnFy0KPII3N7KF0WpmwpdnA4uyyWuMCn2iqhrr94jFfi7VoIu/u/EMLvP
AeNAkdMX6bWvgbiR/gwUkHIGRB9f/MxPCFH81b9agh0B9fW/XLzLfyMstLDD3OBw
vlOn9epHCHocA/liNaXQ++x61oRwdSjZDTEPxjr/uybXZEo69mmrFNFaKXOGr0On
/cslQh/aDFe2HCjt1mE7Te+MIOx5D9UGlaEscgNlt7JPgM52G88PkLckM9rBHBJF
FrtKKtL1Aqsv+H9Vseb5xCRHkY/DfBpSqoHeISYCnMMXE2CadkoR/64AqjKBtY4c
u/xey3h+MXGLW8cFtNg/eF1MFMaq7JvGQ4DOo9T5Wdamcv7s2CULLCR/lo19I8AB
Tmh9DpdOZOkGWil//BlG+AVirqo3sTxce+qUByxLFlpp8PYE6uJrIcl4Si8tFxAG
bWqVMiLVPXhOsL5SQe1Ac/7fyCh+cn2/rQfyK1THa8Z6Saar8CSmUXL4pNWJIaUi
7h2Fhrtp0fg3W5Nc6/Pw8FKfli5liUXMhXrntwSXREySA2VeNSGD31ayXx2xlvA6
HSS9zVT3JF/hNUc2I+TzgV9L7GTwgtR8dnv4r13eDORZvtbxjipZbB+VQrSyQc0m
sziUS8H6wejEaEYeGu9OIJdLuRdOnHmEcw2ohAVyldIB3SreCqbCqn5xfo79nnsy
bMddgUZlXtXpktfw8vSYJCJlwWehhhRTukD/3RRzrQTYhQ1idRoCN7OqIxn1nlAb
NOAR0eC2q0ZYszctUJaYFkS5GokhEknRf54VAltwJ08XoNobXzKgx0ExvfNgMNxn
4k6BOevRWWokvNnHVLrTOhArKRKFYprw0jvyErTIrBLJ1jj099ZeENCUrJ72Vmdq
zt1WE24QerrlJQc8RyAfp3BN7uHtIxdhmcd4nlYI2im2zwN9sjwU83L6PXcUO99a
vbCdDOu1elt94j96tmOQ53G8jmaJ6JE30n/RzfFrs73JDWW9jMpp6ZSDQqXzbR4b
oNeap++MRXmW/W1kq6W28G9JemnPNERIX7cGjSfCYsIf6paN7aFjb+2xvVGhHgaN
uPr84HfIJlgNJnqHO8dEgJ35TyaisngPItZgBKDJZXD5SBx5ZNmqobuzkrO5Ln97
DvMvXU1MwbzsyYe25TgjBbuAwiPQMsLASKVItxGTII1L5b5j2yaEuTg8VmVwe0Nh
io8XTzBhkU2dK7WtWnmgVsUhBech+p9p+BI9c+qBZwQGDvkqpiQifUdLhuw0FHcV
9fKcYJ8WGEHGkoRoNcCUKep0VKWbCjenumjH7Z2SK+dK4l4Ak0lpzWg/zd9jEGyx
F5gRaPxWgqUaWl/aDTHBHt3LFjQwkBcgDFQWMVyXa/XWlvS6N55f1dOZVd2+WjOh
toLJAOZ4Gl3cbVd4WM4fQJilZlom1dG2fYksF7qhcV9LY9HE8vVqf4LQHeykqPOR
PcVJK8WCSyXluZ8jmhmYSb+XFW+2QBcYYjOP0YrrQp9cjrMInBPqKkYLTKGCczky
FhrSBB7xUxdJdhdf3yxfdrlZ3MgKWuC70CD9sSvjS7/kKnM/5ScVwOT6gH/BIwNh
JiKLlK5IfI14/spNzXL3y69tvRtIrpw5y6CPp2ANRlwuqte/9iCmAsGIGAiZR4f8
NuKl9JLNEy2ZLK+8Gj6grOpSqrucErog4/OcVH74JG8bChSxttFPu5VP0nZqlS7h
EkPmd7M1Z72nhtODJmTGBhapSGC02b7gQ4AJxBiZBR6Iu1EGaJx1F7dD2I1A9Xwg
/FxwNtgoi1JO3cPG3DNh2t2LyqEhtYrEEmYfN3bYTJ/AjRD0up2QqgdwgGuDLsWC
iMpM9E9h3qsPBhX07HR+DKKbaNh8QcfPt5wPjHgC2PLgEGN3aj5Wm++5IlCQBSjT
H53xF+poteJoubiRibPEhD52weJiJBL1oP9zQbdUIpXXov6Xh/m3fG7RoRe4+aVA
RZZNDJDQphxkmkzenRd5T1J7RgLYQ+HJqQUoTVqWbpEa8TaqHNWgkMxqFAuPaj4x
tpF20CjsE1GcH3QqVVTp+VKNYtm2mqEyjgMdDvcaEQmb3cLQa7Qu7pUbwbY27i//
GKwHqQAl4DlvdBqE/OCfKAI5VD1MFrwdMWbr3C2LyCUrseiv1/jG8ROAsuKGaEQW
c772npvoIkSFjq6/FO73ZAsiC5KBJHAicyU1UAEsZ+Dy9mCXDymWyJgQOkCYctJL
DmLQEZNgbET52a1sqZd92jdcgcujrnuzU+l3yMWmuveRdEt822vbrfutkeZ5/BKl
UnOuVX6Wve+rbQR+u5yW0DCf/hd9/HavRKOBHEo3xv/3KwXgbbrPxYTUMuCn8hSn
Ow7BrN5pHKlbJnyXOmwnOp5BxU1x+jdmUUJDzagPArkfDlWxmrkbA6Q7LyZeqbAo
tkHx0VhlU9EFxLiMBvFZpRqSnMaOxnv0CgFL0SvSwCzt1wUvEXBBFvCw+nWGfPbO
kWLB4jbIrhAvCktBWPWPREK+ocyRcbfcyN0hOg3BpfX610Fzo6Od3Kmu6HQAZt+R
Jvq4s2UEiiuWSLB6NlpxRrXcv0pU33/kJoWHeLuLiLDKn7jZ3bPrKm+B30gfU7eP
1bgx1P7lSSHUfVA8QXOZIBNsOXWCo3TtqWYxtjTI+P/mI2urLj1TE5ZKV0VwpUGr
ggLommLCleRx6cMTndnOLz0WNMkupilRp2a9bxC3xTkJwKlJMft52tE/ULn58nve
/ooYBLZH7dxARam0eCU78ImQUMwDfjZR8v+P0DfJF8ony1X45tJhwKbOC9MMaX6L
OCiWNlfkllD7Owa1kQf1ZoEGZSI6tN8l9eAKI8jjTiWVglcV7z75m5847o58UNu+
DB894dM+W/Zf4CV0D3ko7gEmpX7JJPK8UZ/leWsTG50h/tCi7NC59ryaGejsQ8iu
KbW7yoqFyxKfsSzAAeehF+Dj22ihs+lsuNISsVj+qX8jrzTn/fm3b6OZfoJDTlSj
C+9s5OX4e847D1m1oNK4Bi23WPYgoq8od02jOltbCnGOnjlzyBxhWYgZsTqYmHUc
sFWZaWF6sSi5dHiL11C6Ng==
`protect end_protected
