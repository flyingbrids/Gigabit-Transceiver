`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bMVSreAuMjYh2mKyHUQeK5FoAtfvg0auv9zsYiuXkzqC4/op2P+6xi49umfH9zCQ
Uaurk6GyJKo3M4WuVKNh1k2pUZzRbz08lRgcUhBSAadxXTTqRv1v0wYO7JYsriIj
8Z4g+xEmm+V2f3lQpdDbqUEQm/iUdgDY7cBSEk4vP4XHtMDBK8EReqAFA2XMomEZ
riHiJhW/FtUpCY8qeR6MMQlMbeJy1XAnfmRhjAGt4abVZAaHGq1dWZZuAIxvrh1A
fciP9I+HosTWOz5fSZTZocxVn6oWr9ZQ5EGLbjv4BkedUPZDe8yzfCDbWA94fArh
ik05TDyz6xY/vLYofmJLUQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AthNjr+THA8EzFWFeYnhwfNAFlB6CDJKbs9vYSaioWHtIrOmKunPcDMihf2W5wPA
mV38GdUe4f29idkNKz1eAGnohTL8RCcW4Hi/Q2kseUwDF4fxFVGpOxy/dQaKHu0+
qwaMfuH1kX8gBhrbRu41r/SG7AXWczy5eQgLCha/TT4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2848 )
`protect data_block
z34ZbEBqIfudlvGCfnoCqMK8AZf0FNobIVGu8rqTLenzFezgKT3UGD6796T0KkeY
lPcWb3QPaESVIsp95eCeJ50EWTzc5yl8imt4eLJd1f5gQLHdE9Zp7MMIa1WyqTvo
hjABcp7Wto1Czfxc92fV4rVXNW5CLiHhvCp2y6fyO2XrkalrLPxreWe5djuk6x0U
YMoR3LhKqvcx+HIu3p8aaVV+5Xf3uH8E/EpyqaOYbfjSA/w0BwjCvEpqsjkKtfeQ
kZbxKptZltU48TUCKJiJNgdyE0cPgu7rcaks/GBAa/LqgSnuqim/LchQsMH9/mK7
uZ0600cLQRJ6xJ2S6l2e8MNNPDwzo+CXS9wo/qIK75kcWkM8DKZ91wBZ3/Qcb/+Q
w5DI6pMo41YoHHoTRH2s2S5G7VlHJqiZodzk5lCNdhvHipm2oT/fGQ3H6pdubIe+
5cN914e7PVh3vC86I5qOCD9N3S0L8uE9zPejZ0hu6l7lRMMsF2himPaA6GCSqoh6
zFfZuzNPIUenFuYiKvH/jMBkm6//A6QDIe9Pd7yn9ZZwIRzGDNG1wxDntmkpbgBV
7f7JlRt952bogAk02G+dno9Ao7RZdx7KqQZcp3LFlpciH+IHW0hKy91XBfFQxSAq
cG/oVDACWHgvG9O15aBaI1tH8owZ78L8o4Vpa9YOKmgrlPwAWHhr7CjbIA6vIYjN
jUCOH16cSAYdwoGqWz/joWpzPlmLqZUyyjMryyIjRXHNayyo3Tr4B5sgo/M/AdTo
uy0bjQHweeLEjT98XveRo/sw9/yGYgwzc9wfvU4E15f5uqUtAPo40bcSD0zj+h7O
AaqM6XODKy9xWkkeAzrICb4K0mGOpcNruat3q7tvUDd8On+AmyRtL9L4dADxvAwG
UrTpObQSYmdaT/PdGKpLU1uH6LwscTjUgBcJzfe0fIqlsA1mNRk8OV8ECoW2slIE
TuoISf3dKPFYYeU1qoiDK1xtJnfPE8cP96cN5ppI9o9L2DKpnNc2ENYgOQJculGn
HJkwT0DMMHLU51P0j9xVwa0t0ZvpR1JnvaFuokpLPcFXDvKqy/WaQ6W26EQRj0qo
jIp+MIh1JjGjoslk6F/0zzBFEdl/v3PrUQ5ti8drzRJOMj80jsdMFNwK2bRaDz+7
xk4hovQlrJGGzT+9w8kERV58cYZJUs/opCBrzoLN27jUlZOlqjwVXoa71k9QhnnY
GyX7HjCm8v2nAmSh7XJnJQtS1KqYsJnEs/njer7qJle6yOYTKnWSXlMvh/Ro/PqZ
xwjX/pfnJQuRXyCh5amrWOctp/RSujYAjkyRq5Hdq8avXkxlaQwRz9GGeGOgBbGE
KhfsNuUpOIWE7Pu2Aj4AD++2jhsClYV6VL+kuUhnoXICf1bi6JI1cheidjbRcMa4
uEYZ8E1WXjozMFfEBDiZtSq7vzG4D61wkn6VtjQLEJEaBsL9+/3d9qBtucd2R8SY
PPfdOKQw/GFoEztoKP+uj47+N2O+1PcKHIb+hMO/j5tfevfMM/tJABHXl436itQa
I19CQ6U6Au2L9iUXrNuUvYfLhHstue4NKMuO1W9ZZkt7ffs+jkMAa0qLdCZxTYsx
w/JwTLDshC8DulQCwgnI2/xpwEN5rNpE6xUNwTQiiT2RLLEQzW17M9JKSmALsv47
DR42dQVkItiBm1/YR7YoJT+i1DxQSHkku5DlHX0tHcE3OEEj/ZewgE8o31xLQ9zb
QFIC/sw3pS9EfS5esqhCE40kMRWr9W9dLIHTTJFPT9Bc+p1NhKj5FY4iWYQ9DkT1
BZg1zwjOBMlAeLbVTmz4LaJICCW1vBdbQn1NSjxTEx6XFUlkLEObo+WAnvoji8g0
WnVWFZ5SpWzdzEOEVZerywIx10NSPUdVK0WTrSyzkHJrwnSVU2jD8zsCz1vqRe8q
HCMVcgLaFAoHFL6qR5FaRKP1Gi1/PuLm1k2syaxSZpsCimj0ckseixUTD3p2nV4i
UOdYQ5xSv84Yf9z4fCJhJG7pjEh9UDod97UQERWly0k54+6ab4WrrXpXRuY+fQMY
ZgQZvqGD/X1hHNMijbbfPu7Et8jTG549dclhMXrxkYkB5LnR9jjJiVMvs+qde+et
YpLUAVyViZ1Cx3e0podrlqH2s5rMtt7JfAWcLFGTj6aa8ow1lYz4e6mKNpgCBYk+
oJXmcJLYefu2aP6l2XQNu06KWf++tngB4rW5ZOqgTj+MECJGmIXhnUuyK+la9Y9i
inH85hgK1EG+QCym9lGMCNzZDJdJMU5Hm8OrSrAFS7qbgUsScUGOix0sH0O+7Wrc
6R9WwdDNXJ4gMmFZ+LH6ekoSOTmR9SPAI5gAfWftwnsR4gzGkc/dN0WM7kkB1oZs
ipFHcFDDd2Cx8CCZZvtX3SA8B6Pl6Us7RtvtCshqRqzi3SCQkQLOzH7aOKJsj/3h
gPIu/9WCqAG5TjG4xfoyTX/A9G/5RWC1z7zUl5o2oly1WRMvgZZcYxy+osRq46ba
zUPXKk9LcnHb7x+epSDNsE80B/jpwnYP4Lv7HXtinyTcZUCVih+i/oxoPaMxtIkA
mzGQeJsZHbenXqP+CrG+lzvVw5d9uPETgQQ7iFoXYSiUe/vz6crCIUsPrRC/pQuM
9AALwKM0PNQq13c4Vpm+LFQmrjNVv9BzR77UH7xjKw2QYpsI8TjCZR9MI4z6FVL5
NSj6qIoL7Jfow13iEG1ymvnbxOeAtf3ER6YCCiB2s5i25h7o/oJqNyecXuFjf0Zf
ySEUcK1xM8VhjWbzBl9cW8/0wNK+TANz/BmI1+o015GaSzxB0BFFjGEGB1YzOCNp
9uBENF27vaaJFVDHxbLfA2QsZtTgCZ43gBIUZXUUYSmOjpCtiMAk8as1qT55eFcW
GNZvhmL3fBChYREv85gKy4FzNxOvO9A1RocjW3SS09zX8M4MMHgZyI9mSTwpA4yb
RTqRL1nq1pCvkQvL0CWxctpcvGWDmpAik0s3GzT4DTCxBKNZayquroZ6MB6Y6iYh
f1NMiCchCMnbiPgC7pWtYZkHxibWzdHaQtWwDN8D4MWzuUEMpZIlP6KdJy8vu077
w4vQIpG1zsyVOtqUU/Gz3OpIy8Yc/m23pPDZEfIweqAmzKRfwoPQrI5oK4BtevNd
BZZ/CRzBBE/INWOo/UGHXhQkjnFzP5hM4wjN/tA/ZTRz5dOWWxyCXnMUzEJB1bhE
MNcKhtvDOX27ZYfyUSXEblTBzSMm6HmctpnhtV1C3olXwe4EVB93PxyYpmlPiOxc
LzWpItHg4jFY+FR5CU5/RoZWTSN73e3FVdMdPTKj2e6WECZJ4GFAZZaHwLqcBW6K
6TH+T3Ikx4UUNudTUdvjsGNtUEczIOD0nSEpT6rn4rc4m2kiG5J6p6kFMsCC/UBs
rZhERFBvb47PkWWURtHfk+Beg37tBwwk6qNGWBvnP2rRk5avk1FM9RBA5ui67iZ+
LZ9naCXuHAPn+7NueYTHcQhErpRtpKppUXm4OFcpqM+Y4u2k91rgcrtSQC+jUzm5
0uwWgQ/EMdhOoiNlQ2t7FySSPL6EzMv1laA1r8Ri0jILWYGJjhv4OQB9nqZNkIAo
T03KCwxBxs7OE37lpEtA8Ee/JeiJX+3sRXLu+ba394ursQIu2oVjOgaEzhNG5ZXz
KYcWn4Sc2s0I0rw4L/cLPXjrY+fnsbQnXsDUUWy05WxVMFwjACE8YqRSpKfGvJLk
dFiqyRqH7S06+Fv2gsD+EjrjGtf0Jup4xb+udRHVP7pbgQkwy5BJNXGNiTH3jBAV
etgawu3GUjCizfaBQi3fJQ==
`protect end_protected
