`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
JkDjQTxOTGlWXbsobqnOwrvcRGy+zYO2TqQu1PP1VpcqamBR5XhATIhZE0ilT6bg
hoL5B0pdR9P0hD4EDVQn+SuZWlVNu/Bz+VLhi9oz2LfoLdSN2g2TZmMCDPAi9M9N
8ZCfTsi5Z95RdmadWEnkoO1dOixpL0WV5kGTB3J6StEek3fZ8fKcm3lbV76UKj8x
lb2a6AsUuG81A3jbOOOB2j03VWfDyd/9Y1rR3J3n0KAOtDhdm2zYCItggS6gDsfn
ZOPgdXiDGBLHtkHW7+TKWu1r0kLmwNdAa0ryCddia0N0vFY7z+LI+ANFdFFJtmhE
RkPvNQJCBw8jVRc8YU0vZg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
c/5SWrBT9fI6CJI/2SMZtQzYts4qNwMafVyb318kn+Sd1uSz9zV9Pme11FDiSGuK
/USkO0H12E3x9oHftGy9qYyYoNiCYNXUiXfAchvi+tJ5qo1rG1F9nd4bF32WcqoL
PU2/+CyBTiAm7ToACT646X/UwDz7lQAdjkTl35rRqyk=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17136 )
`protect data_block
y3nOKM+0Zx/MNawIrrz/yfZjENu5Q1mkUQj4KhZij/s5uBFYxogZieEOj1rJSjr0
9QLo3Of/CAoMNYJ1md88U1j/l3G3tXjM1WkBeY8PbjDt4E2QbGgORm+OnDTXAPtI
OzjAzPJXmcFQptAjceF+RL7lBF1BAPJReSql8uhDwHyt91KEAbaeGCvaUYfHA10B
3tnU3X3RuoNV3Tb/FMnCalJiaVGfD9V4akeeQuXx6hvuNQXLbs+GXEDU4d+kbjyW
DCSY3CxwhIK/hfuYaDwv3gU3e8+1Egb8ZTWCpT60iVBGg3n2AlhJIcMxavf96GYv
08jRM9NWeTsDwM9XnFfmStOWxSJmYvlfPUBoypcJwn3C7N2/+Fu4vVHOV6Xu4rfN
6egO2PYTlWAV/pVL+1bpFtUbDAYUxrqQ4dYaDtk+e3zy6FT/WubTserpQkFk5hjJ
lpWw1VYt52aixDxhk/Sx3n7PDY6mrU23HQaCBsmSO6an3ZC6n2L4FyPlNlqXp5/V
vpXzCT+cIhBn46ELUdtN/2Bls8BJSC7KmqBUOUByhahnTbI9AuXN79WCiAs+OEiy
PC8KfnsooYGPz8cn3LJH1eSFODZSq6nCOtfDSP2jgV/PXk63u43cGokXMSaJEC/w
Bck5OSitEwYqXF+XMzdHs/DG21HDsDyJssmw8Rk8/zktgDccL9R/ceOqnIlhM3uw
VAX+rD7QZZ23hsT8FHfiXp2awDFXMbS5rxNOwDVhMKwjNeBsJNweRoivmXkMqG8U
ZhU03mfZxk+cG8yeHBFNfyOZOBa7xvqPui4cVbdNmSpD67WRre3DRUPjVw8UsHrx
Qb/pHONE+5AhcaPYpWOQ0mciTO/ylJ8f6F2i0GsAGj4x1OQtPmeOkljkY+559IVK
XhMvj9JA2v5ZNP0BMDW5ICzHxFNR/oPU5NTZAhkRNL0tzZvsL8vAof+WyMmd3ncS
LXcM12sn7+pth/zOXL8WSaEA8VDEPVbfMWLPl3nJI7lFb5tBffTqCP4n6Kp31Yr7
1qtF/WZu5lpm6T02UM/cc8smtJQY0LkpMmP8ScmRATXKPKVjsg68WhH2eEzb5xrT
JQA6KDu2QBhuSBvklSRi68M/Lqg96cupyfcHl9e8xlAov7nF+iCKfrxjOQpjTJ2U
WXhULcnDhseJrwEuytiTovu+Z8mSG1PnDLaqgEErunGZzRBu040ED8vRPNUeDWVZ
TgKd1p+SwFuHG07J2we1VBhUggtrBbiJt6EhZ29b2CTNPx8P3Nuaxt3S9ZTwJr+u
7roLjBNIxbX5Pt6VYjGNauSrScKNHF6wybeImdUd2vlRLWERUullZFeLRopPKHkL
/Lzz93XWtMcWf/kN+MsvQtCrL8phjy71QOzjGb+cqsRgC2hS6W9xz2QVsHBVgxBJ
2GjxwHT7n2tSNsmi8piRoOp0PzFJPy2t0XCoSArIbaoSls74q1EpWFP25eFVKnK1
5Qcp6Y1jrug6u8Wb0XUvPtqQnWJLdus9vx/aMSnZQV+KkqPzc866ZrfD9AoUazam
ygasgMumiyh7IYQEGNlkSUweusaQIpx/UoagDIZF9pSKDdjKuWC9GEOeAtMDnJKu
ljsLXRa/SagxMaivLlYpaqm+tDOruGtJWFrdcrZziKoqPrEDZNwCG3V/+/qCcHKb
/K57PhOwSLVhrt6NF8ArTRJdhmUMhqa0v4DXY29x0b6nn2wK8pEZukbuxcsAnHrU
hTa4+atYWQkUhzRwjDkWYpriiEkAZ7/SxUIQm7T9yO4XlYvsue532lKbZ3phnXzk
mCI8fi5zHlyqHM2JZBpKr58hn+eLtEmO833YHei8XEipNorNHhb/urxZP+v5uEKN
eREXJJVw7n+khQEUwpceIYTK7Yeka+vH+xT8/UFAAi8mrJ5mzUCzUdSUKdvgut1M
K5R5JhaNDVg8Bp2vGADiB2oH5CtYgEX1NjeOseFFjK37cEme3HGX5l/6x0fj7I0P
ztg1CEFO/BvR1X4HjwSC2ZnLJGEetd6v8ewLcSJMqg9yLt2qeAMkRlzCIJ+5YN2T
lsNkt5tmn2CCCwV8D4BU4f/w7PwM0wySlK1CE66H3oQQK6uMZc2E4Ya6SxBpGTfS
Zc+IjYffRvggN7UZ/FMGV/eSy/ZgOb4zwZsjGd5gB/HAQ6ZS9fkKuTpGKEhZSRhd
NDRsF1YeKNrya7A3bYLtreYVUM4761npotEcKN5WgRRsfKxTLjGtbZUNs9S6ZzY8
ditjJ6F7HdmS60WXXkYQK0CVA9SAOEV3MrKR+St/lbjp0F7UgeFF1AzpawZTd7hj
nTvL0dYAmFSj5WPMS/zHjJokW5nGrj25fZ1EVdKTqa24paOXOFv242SPH57CHgPE
6bOOD1SlJZkD2gdX//8JIzxgbpkfkI1Ix90Pi87sM5jw6DaVlMFAdw90G/8miQb+
yQXa+4SMBOU/Vl/+npvMsxuhHlTfkbp+wLSntoTEPJP1s6Bhi7mzxaM82fInRYy/
ZQ5DMTp11X/aCM+P2ru6BVIu4UrzfQHsuLwkpzWyjdm3KnAWMG97AMxrW08ZRUh6
ABI0IFi8KTsiN/dLxpISIUSMSBwq197VdzmzoXRsA0x2UYlOrO//zHjvll/9pbJc
7VtAjhzdssUCIwomttQ7k/nsBJ6xZ+YgkjmjhpnkxEW63pMrXA0/lhR1NpHVXpHJ
0fCAYevdBd1NwSW16ySGuFaDF+DK7sebTO9hO2eH5BC8QOFS7rNz95fpuEs2JC4C
UyeqlPRSf6OIDLscUMz+kct5uw8sCmPn/+k0ulD8t9om+W3x2m7IXsyFKmzolyMP
bvVBFLf4mjrsNVFaRepVHPw5QGRgIuyKKbQip5pGyQFBq+eYAIly7eqnECcKkut7
mJfBriqGkrDGITdvY5FOWWxrBeHubxSBBUBGVHr7ZM6pt0oH3PboOnFzKV22HbXv
Qyb45HnCjkrdZYqrIDLm94jCIcMcfNjn8t8EHLDQkX0H6szvQ9sTN9UfixaJr0av
cCmIDjR9Eixx+PNaOC5KuwfoLcCKsxttaDbRdTo1oorQUf916wigDCxJcyuzqaBG
P2uKWjZAVbQOhOEn2f2+hk0IYLr6ZiLpqm9G3C0UI2Zd0Hf4hY+LeSiHTJA4ZKsE
vFC1EO2Vn8ubHhvu1hatMtVgdkR7aR3d9KvVIMNi8ro9PrwHbC0qqaZUuzbPPOTN
4XgtiojPLu3riA4fNQa+J0oLoCJit0RDiJOcbFGlcx+8wtNA4chJ21sXy/iD7y8l
ED4KHSoqyGw5esOqYYHxL+OwDlehEkLgIg99T6eaGSEyWznE0mEtNp+CSirZVyTx
LUgMdhHn93XlALmRHjffHcEOXH5lh1HZIReBrLiWrtG3hjYQWpjdeRr4EyuIhdPp
Lxq2xLGGMEap5H5E0QWtEnydQAXSkzqV4BJB7PLqW3KgEKMEnuPTM5doYzrgW4bp
4mrTT+KUHuCr9PS/88V3vea7TmXiOPIvywY0AvzxUgSVicCym0bb0iJhz7icP7AN
k+W7l0Gt+CFIOydDzJmlkAWcJolyJm7CZSlUNvLuwP0ZPozDNhkP3afoDnfL6m15
3YxDk+VEDjJJeaBaJ+JPWMcl7+5ACeX3Sflj5DbXubGGT1Hg3ACjXledbItADX46
I22krguDgAzWW1LFYiRT0keiHUnz/iRoJ1UUo9Hcfi61GdwWV/EdWlrh8eqwZJsh
6ygQYjYu5C/UJeqSouCFoOgXdNZfG4+zdgqUxaaFhaEiDM9SmWPIHw2+o2DW737h
EkCyhj1ouW1ADUOLfTesgmisKfx/pugz15icpQm3OKNHlMYNSnWjNb/GEvrACbY3
i1ntorb5KfgBN4Bf9FvWR0gBKHtYi7ERbDHppEs6vXgZks4wtciyc5k8qg+pDKz+
Pa8nyZRgWYI7qX7rIVAOPrzAcd11FrTA4ukcRG4fr8dLt/bqSQq02D+JesDafm9m
xzHlc4m3OybDLw07FLLjLvrP9FtcQyztRVky0tnkgVT6lUaQncDy6ckM3z5GKJx9
xG1RygpiaqF6aR+s45verM8iqwNEyopumO+8J2imgWWHpnnLS8W8icBlAB3Idy0c
d6+Pt0O8PYiBu2N9xQ2lclqigPeHaEhro6Qk8yo5U/GKdXIXmh14vymPGBdLOOvX
UJe1weM+6hfMf+QZ/4vgIifPII3M6mmIC6FGJlmzatD3I5ZVnLUY8ICIH0oSkkdF
QXpcZiKzq/WRxNLF7nG912EWGdYcmJuNbvIzUm3iOTn2igIRPX1O+3wpgXvguuMe
89XbkCzAlCqic/kSGSp28U2YXvAkfCNAd8CLl/L/P0IfqzFgqr0qvlIxsPZU7Hmb
m2YzIShFo1dhq3lMeV1AoOjF265NkrosUzzs5H1owkK+PjtuqXbPLk4uPImZrmsy
hQC7hWFrBB/a7lN4slBSBuDhL59vzbQUnQECz29/ymxAGHfX/973ZWryyaHyygm5
DA1v1PBUKVRk9kTlwTiHG6kJAAQpboX3b6gW8dZsrzNVwtpg+AjfBFKHxt7GbMi1
oPK+HWk+67fTtEZLlTsMVC5qDUpLaaRsZHXUIak2ou6o8BHk8vtIPkHPBvDZFtgj
PI+vyV0OGpbuX3JzzOdsbqRvyBj8beoibZgdxWv280jwQmNmHi6wL5vJPGudGlCx
ouhOiyALGzJu5r0eHRQP1Uf4vJXfudICfUMXXTnHtydTReMbyAiUf6/85hb54ise
xDvO9dUXO22r4fbHz72YHgUkmM0yDDrAANhIgv4wa45qda+IpLe/r+Zs2OHJHgK6
ejjIQqSE+XGqafhak22gy+3JUUPSakZtXRFFoKB7VLW3rwPpH3lQ/rpBflkCb4pf
zdjSP0ukV4kr/bmQlWw9LzpJjVJVJUF74BWpy9mP6KOKA4QqAl70qIdoZqTNvNxa
sXp7DQOGpzS2GM5w+bQwgpW4yWFqLdRIMPm1xfWiNouNI4Bdi/GJEKLCRLXJJumC
snvDIPwilV2SmYxB6CrGEAsAIdTYCwCANPi1Y8SZX9Kb8c6zxJu9Jly+yTSbNKfX
kFzHTGZ1pAlwXeEYYQsRoFCfm8R1gXImO0Tk+uhI6bK+EROvZr4E1cSwYWTeGfS4
FR5ZkGX20fcG4kQQeZR9M82myvrgsGjMqu0oG0jk6O8D6WeieQr1sabvgCa5YYNm
QGXMC9oATCdlYMBqPBXFY0BP0USPirjt9Yj4Iyvypum5TlKaw60ZMJLG1RxVp43s
JaPY0iMwgpDGkQklPA4SLfavjWslG9asn4rOQP1PjeppxO4cUFhNXxVl4P1oDoPj
aypidzij8H7TGsEc918R6Y4/54zCK/sDa/UMF2MXGCSOxph3kSc35GDVVEm6aXSf
5hLb0F15W42QcDNh+Nb5RKCko9L1a2TdUNmYv3qxeasjVK3GW4kUzlIM8qCQS2Qb
DNYvMtlV7+XPpIDalfwHGddf4MwoUOguIRyhWiS3FZN24he7HX7VdcPinVJuCjU6
B7KO/uQTdOna2oFmmPSW0i2t0g8m4sQoDfjcJYMZkYTwGFGnb//LPJC5gSQu0Grg
XP/C74/j560nGUj1z3zYC2cW5wkkp/iDwXBCyBhaUFISuVbs4N0H1M31cwKkcaJT
nEm4FDHUmOOfI7Vku/0nFBqf26Q6LtMcmR/cPx/iDeDvemwDfWyjxQA4B/+dlYuB
ga+pFZRfcYnq9msIRMsiV1zsacVMH38holP2cYMvffvrfNNkBSasiN/+Dumwb50m
VqZA5ojf4Gvo08SY69tNPl4cnoP41zLf5/+wwjC/CuDqqsGKh3fAxi9l8JiUNnjj
9QGoawqvdhCrnVALWKBrh7n+e2E+DxjUH3CSMUhbKZUDEsdPFViHQ+kCV/qU97Gq
Tn43cntwHaLCBLU9iYR8ylgMkJQOrson29jEp3IhcwkizRDXYjmgDDjXkvzTWi7S
1YzUIsSWrzhgP4OLCLbojLJKKpuPOW04F8Vubi4qwHsMB4gRK70h9nu1aL27wSzL
b7deOyq9A9Oigekx04EiIiEDS3V8HcnmlbC8skvQHx+hDBpH/mSv6FWINm3jDew9
iBxmCx98f1zlFQ3FeUkG0MhWbGCbEkqiNySFVnBzJfNg/IYO5qnabTEWu7+wJAwK
+MLX0k/2SXJ3Cm/aOeU/u6D7zTFVT28dzppuaQBAyO15d8x/kpkzCwJVs/4/MGgq
agBD99Z+byz2XdUa51OM3deDTxXn6/9B/ey6xevx5iJxZw+kKwXLOeNERZILHZ74
pof+MkIhgsZ/HXfajxbjI5nT9A2k778DkmSial0SdqHJhNn2HwmnWH51556qiMJ9
uy8mYJx4p/REC5CqBQx0mogiklLBT0+rPh+sj9co+cgaVvO8eOTBGO1qXiU1ZizW
iBjVD5PRagxRhVNuI6wxuaE4PXXMENzOSspvHJSHzrgC64qZyfyUUUtNdAFTXwzv
+XqvdFPf/LNxcvxZYlsSA85sq3V3/Zxx9aStrgLyARgDQ4LFJL8aDHRUf4O7jEjx
2o7aLZ5WPeAvSpV4m34w7iCFihG+1xZtPSsE1rb+pXSRyArhNCfp8MJnND8zel9A
Pf6G2LY0xDzz8YQTI6XcyceiP0ytrNXnO3PvZQSsN5yH2Kem1+HGNIOLbseDMWcp
NedMSECaIKGo6xPxFCdiC8m/XYw9XGMAz5xRfV0eyxzt43NIZZV+f5hUXWPuZ+bA
LP40Io2A2b/8JEm73n02Q9CTFNYzO1FcYooUvd4bj/pt+dgUfsbqYRI0CLbzyt4N
o9SrZ02+d9fljLuPo5Y4bIWSXdYc2P0O30lo1SDDe1z3mzA3+le9cJIhxDye7M0G
kDIustQ76OO2ViTWVAXYtOZHyxz4q2ylPl0vea6Ri19/LPjGVNlFj4tHsJUnTa1E
XJ98BHRv6WO6DWR1IJBFfCA6nPGgj/6qyUSLpSh81aoQFpRm1bVzhR65i15BrNEB
WBtUgFPn3oI/ECSsMymDIhsgbNEI3zDr2OCiq1pTQH9fD5ceW2UhvOyyWxxZxe39
QoM69MMOqUwIclCobYi0DrQXk0VwyIEiaMV45urJu4Fo4qdYr9irrMVSxPTcchuR
7d5EWx82qOLJtYoPKc1f6Yesr2VhZ6rdpMxdwqz7GSJGZ6hGkUcNAokiOqA3pzPr
XnK2bUC7qfe1ROjWWdv9uSBrKEn0gl3806WYd2usZ+WWL32RKkVIZjZ7gByYXm6O
Zv8vBGL4IfBdAefj5hbl7gpFqf03fjqOBjbeBM6E9vmBnoiaVe6/q2zATXDjtNeV
K/dK4GLvM+43/KJJ3QIaOB49kYyepNdmek4HP9GEnQSz99GELkcJDLQNa7tNheU5
a6CJt2vD0s1uhKgyeAKWBwNv0D/B6aNoRU5fVdNzm9xITgFDKRQIC/wmr4+s3UsQ
8WfujriePElnJ0O01ep3YDHCj8++uH5q8pLZ+SCC6Ew7g+vlsWKGb4HdV2pfEcSf
9NAYnarDhNI0ytpbmsfsm8uBo/H/xRrb5ZQp94hyveAiweDs99x8FSSgxNjDBLya
L03pW0DIW2s6kjcZ6WDSrU3UMQPfAfsnotlOtuftlqwLXFd30XxEc0Zm3jXmu0bU
FerP7DVheHmLCfkco9hovw6FJS0rZT70uhgFJYz4m0NQICGjBHrH9AVmfspQRuL2
9BdTGKjAmRJp2QfnVPj/K0TZqCIz+ZFjtvrY7vhS1KB5RZiyPjwtdXER1PcedauL
Xxa9UQqgE6E3viiW2W9DLXGS4VU5dh2Sx3ClKnEAe+DGIOmIbhUz2FIn2DfpesuU
g+FxAdIgMybUkf6inc9bOHx3BbE9GmCGPLKMum5qdS/BAE63vb4DRDAKXvb/YvbH
OxhvCeNMIwgSkzcc6mIx2K3bo4AiyEadmbYkXWWz9q3LJug1f86SY5mZsUfyB5jr
j0sAMB3FKgMq+OqIB/Y+F0HdnjlwE3HNp5EL2KcPRxwfN/LwCbnbVv09lO3Nh5fM
6XSfbmC3HjMXAhnw9Oebbl9dpWSlf1U6TGhCvQLyS++0IvX50n0drTMIqTUBVh9G
Se0I70fz+WSuIF4ID3PlnInEFFpQapMH+6YCbE6gHtZOT6QMjcqe+Wj7ER5CculP
13YlRpHwIewf4cAWNH2qXhWhRp3cX+3EPg9ljcXXyTIAdPPdXrjva/MTj9XT2T4X
rzZdMkG1k4VKG58UYMOzsMA/Ba5PiLgnhMcZSrQBKJvLCX+6ttCShYK+cvPBafk4
y4ZTmROvoZT92g7Un05F9sSP8mnENPRQd9P+c4LATrGEPd0MZXM5/Kb9cfbds279
vFt/z2r1Dyd4IjX/LvGIboNRnbTlAZZjjX8n/zu2lT11vpkcvNLWOtz8UawMPA9c
RkJfQGZJMtzB3Psv2rLe/jV8XppoP2EiCCTtot1WfwtyHRT6FkiS1BQT6kH1y8i1
utSqEbHC1JHL+GZdwFjlqNqDEYf9TWua8rg3aW2bq2UaYUoqBEWlkK0TzbEOflW7
u8wo6CH1Wx6XqCxdn3YAc27qgyiwp5hwkmmynhk8QIuBpMSCEkzPUU05KQFfH36/
4H3Yd8R94LuzxPHJNYItF0HHjxWGvRpRM2ILW7a/S1oCpjKbQ0omGZXyjmMEZvLi
HGTwhPzxunOLHuHtZopEXmyumrPDbD7Te7VwkHxLkpmbGIEs5uDi6gO0uvUfv2wI
qJwYjvhPBbiJh3Xadb+PK8nbU4UvrnbZlMCkRz8X5zOcdf0qSPdKZcS6bmp6Eg8C
efJgZVoT9inYOp2NWj3urgMz2i9vv5vs1LYqQRUBKhsrmUvkleH4qioeZG1/2VD0
fqPoik3R31Bs23FynlZDfFrKb23FGcYtHhhSBfC2XKt3InvBrkyjZNqk7EjCMoZR
aZtDKOezcENdVOJFQ6GXCuuu5k6BOG5V91m4prmeTyfGl/RTrLivZbJch+o/Xr21
4hJW0k11hIXwVQNiKJOtCZm9E+hRQMwhHf8Kt7VgXrv+pt0N15ZVk4kkrfXvCzEy
y8KdYZJLlPYXAS2DfwS9e1WzOSwN5sXw+ylerRBF5RqD5F8mD6IPBLA4pY7ZMvpq
Jj2LtKO6wHGNegdLCRoGqDJFJunU2m7aaKgv2G9EdobjazkamEskx4n9WrbQf7/O
LGX3BrpXQn4rYIsiDRPTEzm+FtyOr/KRlQFDUz9jvilHUPNhVibs+wr3MK0lkv7N
wByLWwJdDp/atq2HR487ajF/PhNYa4Cw6jEJkvCe2hggoyEIQkMPIW1d9h7oTtQD
qWPWl3BjDvtQJe42v+qdRS5EvAsyUP7JG9F8Wial2EemFGXYTC/y0kUNXNur3a+h
wL/j2KYSn2mwfLIJjG8PbwmL8Q5CmYaincFk+e06bOFiDg6YHEw67JXMeP+yROSL
YuE4deI48bvuJl2MOIKFahcvMu04ADwi4KfSsMGtKofH1YJZF+rbkSjzDAptKcSR
QK9apuzlmnF3fAufdGMxNE5t0L50RFgZ1On09Z4wNaXiNI6qYtkVb8P4wWnGrhKA
GKcdJr96Ll0xhgVpUjTDhEHlkrUGDI2m0oApvK/fYOfTFjfr1TDsBp7iePrBnto6
C/dnNxyCrE0VsmlEsncGyGNl0vs2AnoLQUfPK1JlJle8lRsElgfsLFft2KcHaqih
FdTQ5oN8N1o/HntzMxBIAbKo8g3F6MhvPFJTirA6PJWqYkfQG83nFJa/DPHmSZcr
X63T5i741aynTLgKOXl3zDMQz9IkdYzX9mMy5hnWEFXSh2Hj7PjCy20kLIaFm9/Z
xJQ2XsOLs8qKC/RhhzuSbd4OXYKa6KarAhLVh+ExAJGu9xjr4L+LfZ+1dQGx8yLs
GtpRxII7pAqUmqIKVLXnJlgPFGypI70OPBC63OuERnvrfR5Fdj6Sfg1+dp9fECPb
Rvyxp7v8fk6ds6miXTRPU4wmKsRPgox7hg9Pvwa402QIRowVzLyyHRHvaK1Irkar
2bwktCjZu6WnAkCwIUHYuwqCucEcgu6YyzdJv6Kvm4G2UP+HtlrKHnUmYubxZJFM
r0n2fg5LlZtTcbxQb5GmRqSUlbY4BXyP/sI8w610UXJFLVFeXgAnSdSUDZt17W0J
x0WKqUXRK/jq0+bj9LMcZbX0LBrd8BO3vTWshabDvf+9qQjHHPGrbI8Exuc93Cyp
GcnOVFFRZHsc1g6ioSIqfg7p4KwMvCa89J8nws4ka9tO+68EYyF9Ru2YM+LTS47x
7aGUHaDc9//UnlF+4WCdKPSs7OHrh519rwj0aI5WF2bmthJMqO1mGMlO2OM9JKI+
1QRihlgjoWDL53sHDCacGdDYueZCpZB8E4Z3Fwed2A/edu3aJ3zUQtM3D/9RSPGk
4IyWvIj6pVeBMinGrkcI9Tp0xX0YKicjD4ApJIfHkxk8ClMx4BELCv0uA22vcy55
Boq3ey2lftI/9fyiVrv1Q2uO98aNKEWZURJq3ftmgpK0ldYQ1LUVvrGv87xxbhGs
yGsLbXn2nwzEPvkix8MBpJ+mOqIzAhnMn3lAyHTzs0e/cONFoEBSP8b/um1ILSdd
hvJadbXIcDZ4W4vh60fD6A5Os9i+lY8x0Fx4YvXBafys/KGSmcvZY+a127GDePXD
XffLRo2zVnG0cIsHiXIbclVia8Wht/eQl3ouzT5BtpYEfjf5BlUbk0DulK+LD/aw
ulQlXO4Yi6cxiLHCXdoJCoH4u+nGHQ/JAplJJbeqFI0R1dANHhidHVsPY9Fr1oTx
b1EsOwEd65tuCduAst7UnxKLnVNVhydDFlG3TvZCoww6HBIvCw1vLKqpl0Xk1uSJ
5RzcG+2gVm09KU1Hjv2lYReWxEMqp4Q2HwCLQW/xSquc3DtGQLD9YxPXNvynesBU
2ASqR5Un/3Xi1kq1jH2EUHHHDtoNNHmyQI5QeVqXYCcehDh03IY0PqhOcp/rO1IH
Jm2kJy8TMgjDQtxw0SvQagCzbAsDltKnwr8zpgv3/QPk+DB2FDw1jG0Gb77CgY4p
dQ9gy9i2koZ7UrIRWmGYivDsnQfOf2kXoMJ5NNyke327AKUbf1K/lNF7Kwccrtgu
+KID2eKdKRT17UrUVwn/vfXk6kwKPcpDxIsvqd1GYt/Ivcpc2thvLVfbmaZwfw+o
POgJFzq5NqBipV9DrhY51e29WYNN2fd1AjoVNcNBBjAmWNlrviNAQhcEQuyxnZXU
3K03lKjouAYyEYfx3Ug18xHFKuYjLGTcRMftLCrBvIUG75Tukk+YQOoAIZMnrZ5C
3Bz0GgAFndoEizR5xv2zB/3jpda/g1PSFak3CqG2V3nIe51JWZjTWePUO/jW0047
pTNdv7wHZxsP3iLsjhZv+/mZYJxLHgHmfUOIJzwWY/6XNmhKgMcSIoRWEUN9rsSI
iO5hy0J3vWHYJHyODgticK1sYV3Gic1yuPOfhAvIudAAfAy1HDjHlyDN5yFHqcRV
lQg9pGCINvbKwukv7G5SD1kGRePd+rmmmc4Yqh74bolYCFRvCP5tzyYqWt9sV19K
kx1nYjWLtSHB+sS9+g7e1EvubhbOH9p2ROBOlfebEMc2Fm01uZr96wmMvPog6B6j
yXKLiOB/8Wwjz9MlnRa+OyrhthLOv4iB4L4oz32Zb114Dlkz7vO/fhvKmpBcPnxq
oHZG/1m8ZkleiPVE/IbOkvYqNv3ogrMGCs7dtkQEgUNiykRMPiMoYSMA6NNKPNCU
BVrKLHloYNdG6Hs7yDAbXzoUXccytuHkJRx3sJ5TOK0jU1f1j9dvm2WWmTBFPZ1R
9UTzqKj7C0NNJFOecHoDBhDxCs2UqLYzfPCACL2cBCKap/Wywht2UAwbHTbMr7FE
5SmRQkMHzk58R+d52EJpNJeqE2RlITtzW6fuU9W53JW/SEtgT4nB895IfduyJtlY
y6vy+aV/IHTAbqlr5yrV0lTkn81pCRiP/EPorbnVXCORnT6OgGv0YZOsk1k7QALO
ltKkPrvTdUy25hEvy8GD/jehrhBHt3TyB0M/Y0AtjVRTHorZDgA5Lt8kTUEWLSaM
SsudB0I2imjSD4L1kAyQckig1r5F4OY1gRr3cHhd8H0mbamBpzgz/Oqg/Ja6Qsnw
Yk/PgstlKl21EtMlMnSFdKHY3aQ5vbsgMAwdQ/WXAxxHVOBn+PuGjV5mIOw+XuPr
7z8FFxn8JlpcGBYeIErSSaYUIVwCOtHerlTbNO175BXqH4gtN42armSsDY8tkoqw
tuLAYtEFKK0MOUOV/3rOQrvdfQbbepVmV0j0PfWowg57qkCj5gq7V1NrIbTZToyl
iZqO6OSm4u53IkH6/y4POM/jeFa3+nUUxzYL6/yhZ0RKIx/UI5/tdV9R1irDUzCP
Zb/pUSA+mjajhz4EMAYGZUvWYjnDDLJ1f0rpC8nPHmgpPqdEvi2PiWobWPpZJzP2
t9UJUATqbQc8DgNiC7SPs3ejBIk5g4yDc0b4nc+eCdo41AGuTCsAxKWQCNIgN+Jg
UW3kR0Kdi3RuC4EMMw+vezI066G+FE+pqrfH6OGSxMlhqA/aNKKrLnwOonUUws1f
z2slYqGU8uap81dRclIFC0XnYIygzCmcWHf1oPmnaZaj27TUKwI1KfTZTuj2fgUV
gGlRg93QfdbMmwfuggeBgJssWBEz+nm13j+dhsY1e+ZBuh9ylrSNfSVLXNjQKjC6
OmOTZ6hB+Ra/rEhBeDoi0TqgO5BwUGkKaD1EirGW0HkjMC7atrhFxCVjoD++WKWZ
tNHxipOmkSO+rn+oJXdVH1SqWOJIMUQrAyQKnuI695q9Gu0RCOHbhtJ08dt/wlLX
RHldN5AvoRAAZGqB24BsMCS2Ttb6PLRSbPxZvVIsHyhVawUWeEBmz68SdVv6sJSz
1zHID9+lH8W5ROtxQAcXd0poeN5IXYHDLxaj9sjLyJl3spS+S2Qaut0w9COEGmvt
k7Ec9VMYZaqKc6dfUgEjkTe7vZl+eu3T4y/osrL7v8GeqgwluzLqy28GSon/XaGO
/DEVrMSExELhMvNzQS1Wn9ffNquwjK+y+NpuDW79ZxW4whFdeaC5bckL4swCkiUB
Txp1mvFEjHBdr6oEbSJJpOtaIlQFFu2M3VZNmODuhNDgpAay6Y3XnTPtqesSEvtA
X47x4duCyGOJ/4nawa2B0udZxpuU15R8/Ym8GYKI7zER3oyo69xlkXQqPNk7y4Du
lceC+8nwlbMWT5x8aHUKU2UUAV3xZCMeK3cWAFEfBRATle+2oCtD7kpbFyNY7JUJ
u1ziNqd7912PFsz6iEv36442/A1tdhaSBB0abzcV1EqBqYwccbEQOJIPciHaEey3
dCcYYnViq8FotIwaS5JB7+L4ABHcmwEraqNm7FwQivCMbIOQ0Aubj4NQd7/H3kB2
2ZcuJYDOD1zGYG4+/Ql0RrwByY/jp1eym9TffjxEPx+Mx2K/InjvL+4G0MgZyoHu
TfWjUBx3rcQzBgr36xyiwy/gR+BcA6WS+IxTrUc3wMnnkYdhCMt8whfhmgk+RJIx
aV+Ut+jx333UwDYX4ZNUfVYEAa1tBFtpgpaMrFbs7js6FmqakiCOR7dQ0UQICIjp
EK8mgA5OQkO7vsg8fBUV92m0F4D5xgDXnZugL7eOZa6wf5SC7aurW12XR25V5Sw8
f3N/g5m9va5NEq+7UiZUg1pmFno4bi4hu0ZJ2FS6D5lYrWaCD6+8B6Y1yPiA91VH
A9lBZcF3pUOuKRgpOBcrIuxWfLcYO2x9tgdJW+3jHzs2y2notT6aaT+CaOqURQ8y
TvaFMaY9lnQRMrIbMqlvoyBEWd75wwfwnVmzKmy8jifH2c2Eh9mtnURuj70c1DJy
wvmRdMbZ5uR1zjRrumm1qj2b2pWqTHIUh1GDeaZSQ/+UcHGUzlWv83YO1CSmTjx7
AsPRsVTTUB1vmejyh8v709rXQe0VCaKXqmLu0cD3aBLGyiyFeANJvon6h3N5DULz
yD6fyulTeHF0zNZb42SWleKzmytCcehBOX2BWSD5KWHVL5VJ0qy5yApNJoE4AafL
SFAg0LT5fYl5xU48elXGwQbM/uHm4VIdXwTghxm5StTn41EFC3aoGgmGv9/rn3eH
nxW56B87Ijwr87W2f+OrbKZ763by+euFpEM/Ad+so3kLFbgi4TaWBN+ADsOArKNq
9+QhrTbX3TGqwUZ2HhDcl6ECC8CuOJkY0guejl/6WlwMjYSojL0iy9B2hUM2fLRA
FkBMVi+2IJ4aoEz7rhN1EI562Pi9Az7BQM7yHg7aFb7iT/zzfwKfVPEXSXYAuk17
dhxNV00gScGRTzEOTCJnSlSPtN1GSgdcuszdiEOxSKm2S26lbsunfuiecJH24eo8
EucPcXLhW8xvOMephGbWQRnkDYlNHflSa5NFe6s8ZlCIlXkWj85nifaRX4vh4mia
YDMjuDHNXMEAlYxsfaKO5HgAkw9aME90d3D9I2B411vKfGxpRzg06WX1xXTDORjE
BbTnZuBOtf8TIxjgJb/3xUgyszJLWUeJgAfChHXpi2TBK5G1Dt0HBBaXzNgbyHC1
pldmIH0ISLZ+1GSTcqYCKKXRSofkClsjmO8fPiM4i4yQbzvLnzCX00pu0oRywgI+
gdWby3vw8dbha31JqxlD9slv7ZJDwxKvHXExF1se7EvQ6ieHY9E2CAq9mb+SQnRR
ZA5fsRVfOlVZZxSv7iFG1LsUjx6ynGmIPzb7gOrEJxMQO45BxMGiCzAjqupb9LuF
Rvb3t/RdtPtqRB6Pt6FF3lfJXiuMEfSMkFQm8MlhnJRMl0nOGvjijaLEn9feVr2f
mk3WNC+7BEZJ7g0CT6nMCjcYOaxGN3OyONk1Gi0gce/qONp+HnBS+vSKBzbyFav7
KGqMLFV0dhpFhxPHoihvFj92kEwlZMumV/oH73KggoOREFu9GdI9nDLq0gXd3On4
rt6/l3hcEfQ0PupOXniNnuOTDJ1o2tlmCdN9eJZ9XhMLgfLvnsGSTdwo6ZXeA2Yi
mzVX8w+CqbnTHCEfvCYiGsiu4LomO7YNcCSuLamnwFwQrbBP7QDl/lzW/vEZnUBj
G7M9GP1K5CK+neM3oCZ8/mThpEwerN8dyTD+LqZTLU7sh6PG+J/41Cfu459N/sF1
Vz7gRRHnj/ojLFT1ABJwFcjld6mgctxX85J+8jfuxJyechLoAgJE8z5afKBVv0jo
+6QPVEI0RFkZbbP5zVWIPI/9c6KZoG38rx9tpQn0rU3mSM/njU1G18q2ucsxhzTe
shPeBjd5HJRXPvxxYCMF6H2e442vrN0xRVQntoNvF3Dzd/olhqISIkWiH91ppa96
toShN+yRdsz0zybkwF/DcDiANLy444XC/22QVkZ+7TEIlc9o/rm1GAuYmwUj2rB+
ngl5xADkPApmHfGNRDcEieJSAw0EIt2tFf8DaWoR4sc5BbeuY5ejam4iP9xdH7e5
fI/3UA+v6Q+38IJm+IQhYHsehroF2Pag/6W8RzKM84Jffm14Izpt70DUvn0gG+d3
NhdJ+BmuvvQq/65lxP4rsL2g5PtHmUgpOYlQgXGwgAdVeN8ltDupB6icnAS//Ss/
bfVR2nyQxpISP29naioRCGZgOw5Cke2Nj8k7INXB15rFaX68U1tKYadGVhnfVVm4
Y2gE0UX9Y+WUKwb2JKgK7b6h22aVFOZb3J+f6QL0EeJc/jiIGNXSgQQ7N3ss23aT
p64dX0j+XKcA1ld+cSJ/JC8GeE1ZeZVvTkgnfxU00WJ6WQZ5NKfvTP12h40K6ocM
Ve1lZa01mnTpeOt6tnDmm8bP8Cg4pJPkbH/UyW4cRIpv1uwjI0rHV5TkTeGt5JkO
gqgyOUyKAsNDMD14CfaZ6UTDBficjOeRFu0fo0d76IDZGFoawIN5fkRXo8mA96iM
g77nh3ZN8737QM/u5JBgJA3pAQMpzwIHJu5sjNmjUxKgTKnriqXkcOWu8pVGS9qw
8eFh9uy2JdOAkO8sABbyfY3ocU2GJCyBdbcncfQjnfrmIL/MXsbxabdlGF2oAYIO
pnq0/8VYriKL28Y+tHvjrKrTg1phcBQ9WTKtgRqhmSw1sxjKajGvspe6TMtglGvk
f+p7qfkdy94J3qmQIE1sTsT6cgEwO4l9/edhFLpDXLy+wGnwV1Ah2zCS8KlfAgbU
6i2NbR5DXCtEn/I62OZK7taxkNKH9adbpQWt1z5j1rlyo/TkIsqiv9b3lXp5Ladq
9yQiJ6n9J94dXDb2mVE0iambTsr1ecOWgqYyZNQ08V7rd2BMNnRLqubs/RG386r+
7mshmxL8amQ8bqfNJSaGgRxOlzw63luidUSu4CuYEASTM20Y6WgXNMud7ou97j1A
jPMYl+L8ReuLMmnRhZDMBoanUvaklk8kRvMjhSYwhz6pPcuko981RHJz3oMQohWg
8+a+xKbna6SR9YqHXFECEf3cfER4JX9wWboaYPGO81IkvgjJrGhYj2R8O2yFKxY/
ZENZf3UFKsCEauFGx6hqSE3Pcc4GPxmWO01thFJqBnEqtCPGMllPi/yaxymnsVir
GBJDIdBXb0sjRX+WonUPA4fm7peceuW3m2CDbuw7bxtHQQwJkL9MJwl9CLt6Z2SC
MXEvtax1zvNBAtoxA0jpff7w/0w7FJiU1stiLIo1LpgOhYXw/sh1+D6S/+4c6leI
BQrYVAidNB4T5jqqGZmPebCgRM6S3gA8y9gj9HIjXCFm1LsufNkyU7qFv01bQYtm
GbttWGxverOgk9mpTUEEDlWiROV4fsFF7QE/yvr81MOHxXhQeYUu1Rv0ILPjbANP
15Pjw7UeJGxvaXBs4o2pc1uDCvA3fnSqWibOf/2JMf0bDFGH1fe73GpaBxk2FOBE
2Oj+NJH7lL/c0hwdtFrylonCtXd9//q9yajBM1EPbT2waQu4bVwfv/MTnjzw4Pmx
Pyn21dBcisy4jaxtd5XdiQI6rvWO1CerrDWrZJtDMkOy1wHZDC/k69afB7jvwccs
ERPTEqe3e2CMg/aY1sv8LVPy1TWW/FluVjQBEA235ucgWrxj+eDL4OvLZB655+cE
0GN0rhenL40DDCirhCp3eaKhluPs/3pjjBGBBCgjIBRklVFdu8G7X6iuWfFIEeTN
7Y/lyK1feEk/zv8J8tPMd/j4WomKqU3Bpfn6s87YVzZ4dfJ8JLsOYzSMMmuf1jPV
7G0VQ4rKTnzccl6aKw+8XEeZCfBe5ZljLtqHZWH+h2l1h0yrmFpV9rWGTfONTF9r
ti43MpysvmtMkXLvampKS70T9ieQZnxmWNZAkUoYW7UFWIflJ5fSsd9Ry0Y1FWTZ
E3WbW7UOB/3tJ2lAPjfqgwhxXYmAxzykivqCXHIL6j5O+yJi0C4Dn8sFKm1i8vho
0VF5I3Of9++haaTNwxM7Ou8YZqjws1vrpbTawI5Mqnb5WKvutW8nkYvPUAin5bjs
KtqqkADxNfz+YASsiyKexjx7dVPv/l6WBL9LbMJgensthJYTtk54ZNKArZehNfMw
PrR0PFRr/bFILltAPdrrp/RE01uFkZV4ty1x7fjrWmlciOxnFVaa4TJWYIFHYszt
GvjHGXk+g5oiXDhn8+PZGfCgfbYeB3as7z1/UjLtkikL9YUMCRMR7S/TPRctAfOA
+JG9BOAbEAkrawYdccIno9e6ctSfMHLzdtgVatWKSGWg60ZYZ9EusnjbqpAIByyc
0BAosX82LbdLfW7eiZVPmnfJRtN/5jhYO5IFnvZnznrPtkEqGsbP1a+3pBinQ1zr
L4UPpReE6JwxA8x74PtB3xWJUULx0u91cbGBNx1P2EA7Zd4+uhmi+cBGfSIE1FZ+
4J7krkM3Pt/PtOj1HUuXX5nsAGI5ezxG/jXdPE/gRwr/4JIpU0ofXT3wS/UYmLHF
4LFB1yN3UhIkyYhvmJSuHYfa/wKTyZGpO4LiDvMb/Gk80K+GVxTsTFNynDZ1ioht
bMAqJcxjE2xS3fPD2/vALd1PK6PYocnJdlx9UttImpTkKGVgtzwqJuQ2OpygY20D
oh6vHDgB8tALyYBXvuOHCCASTFuajn/eWZF4CsGRIxmcO7Ajz3TM11x0lcudYefs
TC+DkNhuJydy0K2MPsiMlsNJ1fTZEpICoS6CgC5LfloKHTfMRyEIysVwDf2Ks2R0
eqJEKdKj3aZ6NJgT4KMafmTXBtya/2GuT3YlU5SHJrrAu0t/vqTjj1w4qpd1HbQ3
U0VD0DGx+d0l/wxwwp5k8v2aeLMTSiiTy9izTQLTUYvGIhOxa78O8IVAkMnw2166
up9kfR/mOlUR9PDTyZFQ78xegRNfI6oQ4EJ7Z0M674VJ5n42tJQ87InFb7PfOri6
z9zLaiifVaHNKsGaVk7Iz4waVKaUAc+z3A6C0HGOynoqLynz/QFQ84e1WN0oIs7M
pgZleTpMy6dWJavlSXnW9gVJaokcd/GCanMvjr2NJUtmeMdkQt/gHFIMR2f6myz2
cGh3nU+WOHYER46mBUsi2dbUOWgWR8aSgdKGq9uBeMLnhSBsMpJqA7EcztDz4nlY
iIOXVMtM3cFAZhi/e6lvwc86i8p7VLX6DP7vT0ancjKDhOLf7S9cbjZKYN7EbYqw
j1WzsNc9WcHmGuup8r6cvUYs2J5Pf+46clkP9Uyt8BSlX0l+jDmMaRXwa2YKJioj
CYyHjd6LlCTenk63qYuPb3waKWM8CoJPDO2sRBDbITKxrHFTJA/8vnFNXD+UVM61
fG5IcfDBCa+KjaDaVVeUYhwE3Xp5C3NP9jSMIxuZUh4o2/tHyGyzNy003bMXP7c9
HsTN/NK7bGZHJ53almnNSaQyrVpwc8Ovidw60TSCAJ0ECjUqCAuNOnkDmnzmAewb
T1bqnbEgAnPBkoqYn4sm+/yxP6My8eUlvdEhmk5FrvlUz9/cSoDZtwWkTN/G1tNV
6kGiWA9+4w0ORRPy+Rr7u24j2VPmO/XOueLOWF7PDDpFn2z9eSIXsnP7gLBnbs06
QiqFz7FXnRGOs41+4uGRwUkKDyqI6sAG4bRuZKvdiQG+7Ad8XUih+uYEUzvgKiTO
jhrvZuf3waX7knDHnklB0TXhiKN5SLqkA79l95BIrOaoBPO1j1m6d3eqW6fExWM8
tSn7e86Gr6Btey4QaAuW4nz6nauxAmK3cPW82XIIogHbBbCb337yv4KqiT+svbQc
D8T30xN1cwS8UhDEvjhwIGKb2P1+ZuO5mIc+5Ry+5JLOPaiC/bTXMMZkln+vBluV
criJXjuiEE1sFCbbhVYg8t/bMkdXD70dSPPFD2BQKDKcLyeGTEQg7KrlrP/bz2Ry
t2VCwsAAXGUoNVvaCDhoLuGN9Dn6NamEs11dwm1Xko08R2Gkek5fJm9buO5GFKcg
CQlHoVQmd0e02p7lMXijqwZbuLtILMZmU7ku5tobf96KG8bDy439vS9yESzDHflU
etyqflCEFMsggRuXgAUaCeqDtXN2gaGloY6ohgt33AHVtVo/vy/NWck47CFv2jLI
DTpuoUzkxLyRjY3L45N202JEeD0QaEjnDQ5mlfyyn7c7Y7xzzLEaP+z8CKfdMtcc
NHL2yt44JvJ0s1TkP+ev1pUP7yd1gh55a5jP9stTmFVfMDeRBl9WCzGWszVFLZ07
1UuhUYILHOBMU0bs1QMJ6PlADzInVzMOXL0EVvXzdVRbC/LuYFW+UoX70DLySOgu
/HpHQB0j+rO+2c09zPlelNdJ2TFZuEiD3g/hpfHS9IUR6yk3R8M7ZA29X0K1NySi
BJiP7oAnLyelbktV0XXYuCJMSxoGp2JVuwNesNbrSoDLTP8W+ciNYJr526aIGDsX
JsjRVBGjo3hB2LDwUdY2eF8Ock+0G/ICqWSuIpFfph7ONRKFw6H8nTzalev4rDV2
gpCWt/yFCyDf2YghS1oGrVyUguOq25rPjj7wCjbw4LuW4LGjEdhhqRVgvgFxkDpO
4k3tkbPzidVTSILrCpNdFoUbSgAu9aJlaJksu4TJWCMH71vuMJo06rR2aZ3285Dr
yFR+PwBP5S8c9cBYoj0VASv6HPVCIaz+T5LFrR2wA2cWU00ivGRZO9knmgsW/FSV
CZRHkWavZn++LQkEqeAh3uaWNK/QQuSlECOOYjJhrGa5hzqNZs/1jmKHwDX7Vx0+
SFOJySeQccCyQTi2Qx/YiYBkDZFzwqou0Th35WsRl6uiT24hTcRzlpZRoXvTCi3R
Omi5pqgXv/qVLeT5lw2+yu0Q1qu54vHazksSmjtn4pyDoT/njbUkr1f3oEuWawpD
4E2HcxYYH06viU6boe2cpTOcunlNaZOEyZSLN1fhRW8RFArQjp88rfH2z90RESZC
u2Ougs7WIreQw5fbTZ+9Ze7dMN3fRskMgqyZe8mwifUYMSt+3P378dESGwEOFGt3
fkJgD8o/duwATyBElAfa2qnornvOP2dRv1LjSXJv8pk5Kny9RoD407QZ4NPOBx4j
CJmWRkGXGBV/IhmMlHCpRav3dtIuVZ9xR3te9X04R6Fk7V8SgLw2+fwuJuFf33ZF
jbFqFs9GbcW/OAydyLJ+XSO+66txfzOrOPIY4EzMXHH1t+dySrelhH0fCUWqozaJ
LD22hAH6MZQwCVhJY10x+RCahweV9lwIybAVq0o3mzvJJhXMAAsmUPTTV143CHx9
HvfWRbET4oCIgg5o851bil3I/m28OiC5RP1iogWXZfYVOpGBpsT1GrnGghIshFDk
9OjCdiq6nOwHtCFg4kCYsOyCB+tSUiBuULamIpzAHQI6Q3QiQAMuzyAFduwz3hSC
y8hYWBx3iEyE02sEOZnpItpZihEMhpbRoYeK4gOSI0nBkUjBmtv/CIDcar/SIfaz
3H2jWLsJ8hJM/Fje3jteTB1ulsaSGjSsXZqqNEZUKfAIcRK/jypIb1whEYPKMUjH
cm9LABWUmeJKKVbz/0xy245rK3nkfZUSG6jzXqwfy6qnGOUej/qtUoiWT66YnEvq
I7Q3Y3dAkZSI3+XWbgxqh8/BoQl456GTmXtYFyJdkstV5mY+UnSzhmZT1etoJlMk
IK/Dbslo4WhQ9vp8kEEqfIlCpSCb5LPTgxTz05ZWPuHuvs/smQkbylbxOhJsrB0O
E/em4IM80ROxB5DmnKxPmHjYK3lAoUsWYEM4kpTKb0klF5GLCmxoSBt3VQ0iJ9MO
p+qrqdTK+cnSxIT4jLIkgHqzvj9+EN5Yss75uoMsk2ls+dNAGlq5T+qFWo7lTKu6
EQONKHTZoGseD9W9PcciwV5+AK/ze3Y0KeszwurGiQagprlI5kwk9hse8u8WwKsk
rHTWIujhl+eviBO+9OWyWtNHqYC5t4p7cgwFCO0EMiVebpnE2T/C2eIUewHl/TL/
nxtYcGP4JXFLUOydn4FCqxfcPzdDebmTyCt0VHolR8xuCYM01s0aHF5yljuDSxYn
fHea71RnQCipbPxnjOftb1STTFGQsFOe81LnVVhYPaJxXW7Mxkm4Kivg2XMOjKJN
QdpUIhuKvvZ5xZQK/5fLxUjcq5lpv8ZLrpoSukCHqQYZNvzo1353KQr/cegyi6ji
JKgjExogSxPxbbX24AQwqT2Jrb6PpvQ6B2k9G0qRNrlsiZ2CVYAzmV/tFIYJ6uvU
xlbtaCjDZj3EICTYRHcQxqwdmVw+0MpGZ5sCV2YZedUMnOVGhPo78YkNTplqDK/C
Azrsaf6SVSIZ/xHGHXLM0zpdTUVv0dOjM+/ZWSy3MGWJsmEVD5HzAjTtGTp2A9j4
e843B1JaTc9LE9o+s6QnGYFNGCISpRrVD2jtMpnCdQ/rroMKX780LZ6wfiyUFiTy
tBID3xST6lSxkHALfTFni2eGttD4GFdjepI/DicvZt2r6E58eWOSA0yOqBBTBQAF
UIDTmpQIPDmT1a2n2MF9s7VK+IYXU96nU+2mdqnzsb+ql282c30E4tL2OCmex9Vz
02mqGKQO3nu9aFXT67SUspOxkw97yl13QdDt1wEA594lxYm8wm/MsxUSfvvWZKon
TJFObdJl9yYci1CA5ak9ZdWbktOt/LtTvm16w2E7DKKNd5u9rr0C1WAWrr+Iggox
C461/r7iVf+hyzQ4tvChWe4vXiC66tEtbzcc6TO094+N3OZETZmOQ/yIVP17jiq8
PVxj9AgVHxeMB6cGPm0W/PjQslT/Wa65zNpJt2Vc1aoVMgHJDuv/aQTAnjrx9/FV
kzww1TyYIKQ1vS8d6zDiAFU5PTV3obZ0/iKWUUvPpUzdKxk1xVrs36kx3+wjUTEz
N17BlAmaeBLysNkGT6erKham2ejcvcikOs2YzHx/qzS7XvQFD279iHJbOzGTnYpv
OKhq06NmEDHhjitcGgJwNCPZJziAOflKf47gO1OlNGu7MuKTP2HGfZzRAX4nFGlz
u/SfwTU1sgYQoiYW9ZgQ/xSyKE94tfDsFEapcp2HMCVZx+Rg8YmGFN6PqE/eubZY
gbnNFgrwaodHzDp1oO/CCBcNWOx7cnWhjtO+IXvlcTe4+j1SGzVDEgqkUjZV6795
iq+vcocILvOr/JSKBlUxL1n1WcZBCxBrgyY7vqFF1PKKAHz0+qeRslowOh5RtK63
bSyvCYk3N7afWR+0x1LgT31Ay+nTS5IkAvqh2GqdJXRyoAbnbXb9SKhJjiEB1e6D
xkW9I2/GTnH13gc/TOW5DTa3sbd4Eo2f+yJgw7J/lrw4k7Lpo2Keb1smusednb2l
wCeDBclqWA41wTOxfH51S5Lun+oij/2+OTaAnwsdco9xHiliUZIAmFS1vpPkXgSs
8MQNXQvpTH4qjJNy1tBHxKuipeJJUMjplBBhZ6s0R+XgD5omiGkeEhA37G/6VNB6
U/8OmPRMO0Ayc75E3jcMBCp3y0n3pO86RC47w/CyZg0rx6yfkeX8DJl3vonu4Fbm
`protect end_protected
