`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
P0RckFjEVjh9xjEEh3cDe1HskF6PDMnhfgyKU3sH6P9ysEJjvMH8Sas2HanGizKC
2yhCnRCQPyWXKyRtTa87DqAhARD0eIG79L2tkODH/8LcCJr0Lhi+THCkRwtEgU1H
5hVWWZhCoHCDQp76nkr4rDWOg2KkC9onzajNCI/joiItnYczrSMm/7EYKFLlX1o0
dkwkUua3iqJmnoPKHOjtQ918DZTu1bh7wVM8tR+2WEC+0k9c88e95LufbKKpl62s
S6RbKvmxwq/hIemUxXXpuc49Zex9++XjmFb/WVaJz4PHd46WRkvPmkQXHPyK7HyB
TcDsQUPEi4RJAjYGHP8mUw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eW4Knk1vUYMyowrYsiYabpNPXIK/FfYoYdhEjihqJn8eLkDCgCmxU//KlYP4XJCV
9JYsOH+T1+igDj7ngkpXDmHBUQcA0+eiieFwSE2RYJx2j55JoC2lHMrQv0SiYqVs
RWG7S9YVcMvvWptYkOhfsl4GAxoHRSbn4CiPpm8ag2w=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17472 )
`protect data_block
LKvHvLW2tYN7fEhXfXVSqyuAy/IwzJcqPoC7PdYEE/V8epj2tktH7QawDAV55hDD
JMhs8WFyp+qBcUq9JnqaHBrp0W5FJU9itYPzA48mn30M6BNIhq6f+GkZB7PSMenX
NTmuAPo/Ehsqvsx9gtLnHW435M74AGi5jgeejwzPeHLBch8Stdnj4TVvcrc74yj+
sOJ4j/cnWMRTBAwV+6EIndeBpU7ynj185yspJVD3YbLfOW/DhYObOz8lZJFeooJl
oLHRv6bLS7WDz3mtnychYKK4N7ONu8VEdn4xAeemR5+pYLkFb6ioweHpsZOs33r+
q58ffdMohTbRQlgP7Z3IrmATgmBykuAxZxAtQSIKZBi0mHuCiEdOTPwDTu/Cf+6H
ebbQD/Z1osibySWishunhCB2Ak2Mc/D8hFBzcT5AHdlEJp/WWzRjXxBHjIkqQj5P
GLQ5G+Zx8xdpyzqUePW9ISl5PspSGNBen2NDKlqasEVQ4zojTe+9Rfd3BaWHiyd2
T1tkZfHbYs0PnmsHhabZXVXariJ5SCPwRb7+DWQdNp2Jn0HurDEjdZWyGpTDtevi
A+Wc2Gas/qT8aetofmRPbirLyKLirAAMw19xqjc6fmVBLEFxC8gpmxb6jjYP4HHS
Dd3eC1PCNimga56vop6k+2bGh/thl/6ifN7K9tYfUxC02HB6gpGChSnxkJJXmaj8
GGmxLGMgjcPoqwIkm21Ry4HioL5Kp9G2kCJy9ZhgwFAExm9zIblqCMKPjmGTqTE2
kuOiENADdwrvV36EHShzv/CCF6YcYlzJYAsQZE3/iWrUVv7V9c/LybDdaW1eOW+z
L3KueZeGAZjRwSaex0WqS6e438yg87sC0FTp6e0Fj/7LyW1g+HQcNjNmCb1t30IZ
eu93GfDcSXkuWT6IdQDNMDJQjjWiA1obvfPahSFZfPIShLuuiGVayH++xhbFp26r
e/Ef5TLBvpSw5sz1DGoQUvWEg6w/VhfKzRzdrV+1w9o0owBfxHWBcYSIbM9dtaNi
Xtb2ax3KGHjGt0hZmVe6/Bxml2W1myFPYyJUB8hOoMKCNyyMYAAw2cRcRA9cE8OR
pEzeExncBqFJOZ/HyeWk2LhszWnMMVud//WFZ2KNtCCJGz6KVnZypzLsvsW36CZ4
5fNOuWbuvis7nkfyNoChxgqrs9mShT1nMikvcxadD+6cHso/eFRFRXDsTkd52aCL
lV4A3l2yS43QdZdcuN2rbySdVjqY/bdFsqTK/BC6GsTdGVk1L8bxWSt0fJl17ALh
urfV9yR8CBtioamX/tpxnm7k1gW3QEZ7T43YolSabXSx/voQKKjrowuqxDS83tHA
eLTmYA8H2haApSGlv1YguwaHv2c1eJvki10xn2OcXHVYcY+G8/o+JU8fVynPrM+q
JSqCGjV0vqmS1+94XdBdTd9Z6YDhoFS0C0783Y59mg7q2vIa4eMSqhsVr0LOQXgI
/C6FN9jQGouwpylQhePdjkwP1jyH0F/aPrsAf1pM0SQcgcve/qGlA6cSX/zqT3Jc
OgN5Q45oNdYYH+pJZD7Skl834gbBbHKl08gu0wt9md53s8YmFE5D/LSkKiW+WgmK
8c4cgXEybeg8eLQU/S7wVA4mrOIFo4pHW97N2dnqKe0cT81n4Q79bDMQWIjj6ANG
ReQojpx2xPoe92YH8q/FsFyRp615txY5Ip+kcEN3dDB8PV9Alo1E4LKWz3S3oHgf
I+kqxdhWkiv+2xwdXs2Hfct52ZZPrsYDg8nUYqXhaLLhq7dpliwrTE2LrqQHIcfj
JfiPLWRMTJuekuxPmu9mbpxw0e2y/2H4U29dGHso93TqqOyM9M7hWOcI6kJHOFNi
4aOxzRy9vRYoE/zZs5WWNo19EvbTtMs4ay9LRgM3rRo/qmE7Xpc1MH8osIdI3IyZ
8WKVcVKpHzfzjDfFQBGZuNMVjThQi61mnchkL7zYDgKrB0tkU+uVPfvbKZayz394
C55Y1ykItIhTNokVMeQLL6eOp7aGbwJlg+IiM9f4ztFND9LPtAQqXjl5VqWF6j/j
qyckceSIXPrqdjAUyeyXqTmHeoJxC8gMvTXhjlWzL8rCPsazCz6vU3fo+GJeMgRW
0qJahvh/+zB7vwXkHn3Rcu70Cvav9Z4zo98s3sFqPTH0CQUffcg4Z8xJMnasLZzb
yo7kg3mZGmq6xb5bFJHYD4cKCZCOuLOjwmoA0jEb0m9/+WUlsw/+s4sKKt05+AmM
ccHvFtcXulcjewaKn/R08MG9XfUW2Mf8JaRg7vRfbNVZ3zHrxDzXVpwGNIco2fdd
3pHNMXblsLDG1CSMv5f3+mBuAVsYjs1WkpCDoyvWHZVKqfNI4DbcmbZEMOKNF+T3
N+3HUNO2279X6KU8sarfZ+0pHqCIAedEJwsZgvf8o8ZgUFGEf0rDC8Xbs6Mr85eI
n7aPwT6Tmzw8ToYeXDrOCZvzAs67wEL/UkIskhVeBM4AUsUpxVnPnq4vX+cfu1uA
KMVHabWmvpulb+Y9cVgvYBoo7/ci801bQZxBdc58MJi5XJV9ryDTFcXloInLK+kn
oETgioQlVtvdtLikfvxZRyJTAafY7OTOoUNT3fOJ9B2sOdbMHQ5lEtbwpp2M5Zb/
31+jJ8eT/azBl4zNa02+SyFXz1nbAjEEd6EJdPG+fKQkEcw1gJZa+wlA2rma63mH
p+bibuFCOkk8yEgoY7wwQOi0RTOaWgsgrC7xnuxmcMmCwVfbbEMwDgr0P0tESZOy
YadkYSbiwjzKyopOHbWYKHs0bKlxFfQ7EUZyVejkSaNwtkqxet4oWRBI2oo1j9w7
o3rJIArYdVMxlu0JiFquC7WxNMmvgtttmaidMY1/OrBpIa5izLygvHQ7Sj99BW7t
5V5u+Q7lK/CW6Y3gLurzQPylAgIKT7a066F0ueQg864iLBvyo/lWH614VZLxRkYm
oEUOfH391elk/mEwXe+qe0L1gEglDA7CXZQ2FenDwVkElJyBDhaKEpzXTVv06lDi
JBxt+lUGZWBEwVK9iAdr6kwgnlmiwO8Iv2ijRjLkYbvZL+urRa4hELyxPjtMSjb7
7vCJOYVMrmjv5u0AHJpTmMj2QgRBiFoEMbuw2lvlb29J9WNEWtGp4K0d7bYJcg4d
tW0BQGCailk2DcH5/IH44Hp4bPxzW+mBFMEsG7BBYFVrt9Smqs198DkC5ZBUraHW
3bRBnF9fuw/Yo3FF4e5FG0JwWYjFjJH9jPrZMwOwRGwblgaN12dM0+oWuobC8NCe
vt20YM4aznfiaHb5tewXU5en0ySkAvjd0O5LQtI3kuuz0DDxHLAxCnh0dQpYA9yQ
neb3Ui8ue4bUXmD7SpQyk/MhKo+MZfRs53N2O9KKiGoUfcb/TFGrMxYn6ptNUDXS
ef/vC6c9fs0rixZuRNPKqxT+F86hzKR56StwK2FXU+T/WI6RPFpytsqeo2uf7Lsi
Exa9cXmF7IcqEi48IyHhZZ1a5985VwNQEhJ995nyePvFbfeEfP0MOgJyq1ScWh3g
Lx28WuWnwZAUrLNGV5nlZSO9ywl2Tvut/S4qkElWcvjYg8X9O2JxQ10nSV2siG1L
z364BNgyjiVdEi7xBLm5wvMA5kx6/8r1luoAZfKxmMwCCS68/ImUDIXM4CgWmdPj
b3bXQzJInnM7WNbZrVyvIGJjFDiLbTgULB/OfcKtsvcpjXgdEQekIXqDQ7kI92CF
6alwWL+GJur7jIbiI/Pf1Uerwdhb/e97a0LGw9ofcxVSg4DjOJamr4wmAW04FmkU
RlSUaoKJ71uHwa2jYqLA99xiN5kLW0VU6JDooyyagHCPG+Wrxwh9434xceFIIkg5
VsUa3QqXZttJqIvK1EsDP0jW9tQQDZ2lNjCKlNK6v+NnUBId/yHRPybYfFwLLTIL
uLjxhcBLNNYmu/w8yc0V2tpfcxgSTHNSh4+ngrpeRHD30Fa/Vv5j3Bd+nijUrfhX
BuFQGeBttfJGPJATwDdqVWN9yqsLBY1Wk5Gwj8pI91UGyLObmj4PwEb9fsrWI0OJ
XDydGibkBMLtXol1nED2a+OmMNMZHWawSFewaWGrOTLgVyFVkwCA15WbTGhVUlB0
SkkhUcbvAJra8PoFt7ectuM9lQMYxCrUrXJg+VIZ9pEoljMHozqJ1g7/aHaKHze2
ZyZ8BDnqF+b5PedANAnk0MJk0fjUgJcNJjlrClksjAmGGmguOj+XvvFJQunTHfYG
hKNqtqmEAPkHrw/ttN2tGbkBma2zSoKsJrRz2gt4IhrSWKkJVi6AtpIlOEN/zaG+
6lRYHaqN+/y4VUpntN1SScLc7x//GzO7va5//MFASZ42/0ZDjRxhORgg6zeFRG9F
OooY5raIAqm0MbJpOWAaV32szGBIQsgWfZub4rMxwxTfIj6fZD+dZkAWLrmk7K1Y
8IZhxqzIWX8BNiR1VisaL7HpAcaq8KMSKLo4QcGnquYcxP1nK9xYVwtj+a8B2ygz
lT5Y6MBHCaikrVNIB3o9qUoz9DzfZApxWm/ekAf/2NSRiArLSNZ3k9k6bpinJbgh
6KPC3jPt4AXBh7oAfCz1+wdjb7InHIeUlOqtyIWzSBj5mEUAT8diqMY9+9q/k/0A
kgMN1piF4d44XAlyFYq4H+IaQQI5eokMXtg7eY5jbqiLctSbMK8QyzWHdxlP5+TK
bGgm7GnCe9l6Um0/R40FlYAADtsLH4LIOdJTjXnNN6hk88yljavBYFnVpgBIXQBk
v1DRbFpmlI2eMMxu/+sMQTLaaU9UDrZ5/hwNa7On/96cnNAUvakXv3uKDrJhmZ1h
lunMWTV3LnwCxJr9WdWXKcizSuztxQpU/6/c/cBnVbA00Vagyu8F0IZHi+h97F9o
vmUpq1rHAaOhLLJ1DPtoLS5c8LLo4MkLs9/KE06QH0U1XL9RDyL6HZNTlGsYnYSe
UjPdYBHgFmXWVQedCXRaa079+Mt+k040YWiFbjtYmxRdioUKsKpVxaWq1pU+R1Yb
+hQ7rmmG03TySN0Zz8UYiJHMDY03KQVlAG0qDN7Ljcp4XlPQN7hCe4fIpVNTSZ0b
kOUL+PIXJVzeyL3ccEA6WD+M4Os2Rg0NnSVc03nTM18eQ44gOzLX+NFLfO4baXKx
8GfOmMWaEIcq8xYuOCIad5IFNpcWCCZsNHvFbX6zSzLhDvDk7tfiwHI4D/8c3TQP
hSmApKmpv6tICtzIz7PHDxwY/fV6eOzI/sErKakDOKMYe5ClYqyWPFZwyBkFK3+8
KLu747UQoa7NNaEONSA0kIS7b1AlSpkRemUxHx/C3cXug7DW4bC9tNi7hhoqNp55
UUeLCoXgT74BsOd7FaINRcepAGswJX6G1u8m6mkBRR79+DfCXA6FMaiwyeidrEmk
0vW47YPhql7FCYEJJ6OVw4M8RbeNMWZYpAyRSJ+Q9xdWuA1aAbXhBXvhG0xeOook
iyuG1oo9heaSE+1yaetg376iiVJyooSzG2uKlZq2R4GtMtWbn0hyeidW1LR5XMl3
OjeJmZQANvMlBKLkuFpUE7evfiRfa1XaDwEucLl+xf1YUVS007a0y0Xo7vk1ERhH
R5l8GZynwhv+NPle9cT9h0N7S6d8d1otO88GD5uXO7tROcnQJt4wF99ttQAGjyPn
nBNPmfbb0PM8jfCA0KyRYV5B5uM+2ALyUuJaQhq98IhAqhw9UW+NkoPRoGEYnKTp
g+162OoOmVHwwNfXTzuUA9BzLsU8Imxxmrwr5fPFca99RMexNkvMlmyx0dgegaXN
QjI+yTg1d6hL6iXr+/pZH3Ods5Hy2+eff6BMnlO0ClOe8kwWvwSH0T1+D02IK7/z
vmlFmPwSaSa6P0ntnJy6FUO3qUoXfMnzvE6BgpAV+NFxZ3WyfR4p+BpIeQYSTm5O
yXj7c+QVdvsyfa+dGufi6XmU9GHTAEdWlN7etoKHBmBuyINbH062xYvuH7UEwq97
MAd1586l0AlzElfOzj12EPi4Eus7RT458VpKOAF0A0PZQqDhnvHB4quKOQCqvSr/
wMlLxaxGBV6HOXXaBVikyBX0PKjDAzRLAQg7TX+oL3nZ5qSqXJYeBjxTXjjS4d5L
1koaDHPQ/jUSd9t3dNA34QbzhfNM9ksuemqy4JvLOiRrjCbl6hw+DvCrpfcIuFL5
Hfis6tURHalIBCaefHICabT+N4cnO7FEzvtf1AWIVtNuuPTFU8PS/O9GnDKJQOwy
yEe9FDvrrn+nD9x0OjlbuOHKMROGsUpYyGB7qrebAmM2DiF7y9Gj/rsjD0GuyZdU
Cb9v1w5VrsIMraIT1HdDl9aSwAO6tWvSkB9gUorOMgrHk10PeGnDNdEb3EhJNkJp
VbatuvlTdz8JzXudsVbDgDGyhHpl9qV9FLL9gHn2bZegFmt37t4lQklK1Zvff5Uy
jS1C8w+EQejWlFRzi0MNhbCOdo4yuVd/dPI9hbK73TLeuntafadiIURfXdSds7mB
mM6D8b6VKUjvcLq5qVfkKzqN645fppgKFOD2fSDb8goJ9rY3wNu7sAlrdu8UBq7X
riTy6wjVyLxp/Q+TqArKppTTMfTAXoB8+DLM70ZkxCqX7dGG4NNThHqM8q7sF8jT
J/0NDZ9O4kxnp6mhGUIErb9Lvtnm9ZQpyk9m3N5uimRpl66vQR3KaINt3quFGhXb
laAlXHgaGVzycrjgUH5vkIrq9By30Izv2VLeNPTOawGiz/1GxBrkaclEedGgg61v
z5RURKBjoOkammw1T0giXbK07X/v9QTQH1iiPXZVbAAphlRp3j83DSAkjfOvT4Sb
aj4Y5+o0sC0nTMABEgMxEo3PGCwQmazzMciG3b6cnDXh4QkxkprdhqSWP+gh9V5t
ilnZqXmzECiqYM6YVrwE3x9BQORc9U+XoEoFvxhUiOa/XSDh2Po5GwNIfkogNPVu
v3gkGbbptc6ViHSVBl94M72PK6sj0JdMit5qqSQCl++J/CV1Py6unBtl8insveic
BNPqDI4WVYPabiue/hySDvNDIMPXorQhD/WR0Rk8/Wid3Iyu0Ejia266QFuTzpyE
Bi4WjFOoP3oFWm5Ki2jg8579pbzcrTbrkWE1uTwq3gTWxr7qlMsPCKeW7Be0+9g6
+fMoZ0tgtGbal5nRedH0QCRWzBcgu1Y6pJzGJ0dVNX5T6saFQVhbEb/tEkicI+PE
ucsy43uXcZ7FIgquW5I2r2bDIEMAUkr9YxdZySAe0SZv9yF1//h+TegH3n1vVnEh
daGjgyvOP74fuTHNnWsk/jow5nTlYv07jfHMQCnwZFmkbYLsGPvevIjHY1AmhWSm
d1MVzLXw5iGUbRoEkOr6xzM6OlQtojBhyDiXkCW+EM2Ub1BUCRVvDTsTROOHOIaX
TAf4+449gcQ7MNFH7+VRjrlEJIsigSdHSyiXkmDIJIUEKSzdloXVtSXEO+DUNgjc
6C1Opp4sYJr1XIg0mu/xHLdOTykShvv6tGXRg811M9lT70FQEzyXqxFAy02B50o2
ZUGPEyUYp2blsvKkMf7U1hOX8ekjUpyZlbX5ggVa34HXjFM93ErckYYbl6X0QhpY
ooY4WPo9NJNua3FPgyLsI4QRTj6EDPII5rED7hQCnxsukQ4xU1KBpvFu7kmOjsUH
wSMlTXlKvi72qgV/N6IDVCPIw6SjqKNjW4eI0IZnSIEAVXcvORQB21i0WzxWPrq+
qT/LcLr8miQCsG52eHL+avDqlKL30LJFh7aeeEk9Oqwq7BEJO7F0SC4zZgDnQ/Wv
DXlMbq+zgEqXI2YNbV5u/Q4H3kLiiwbLeJ69cdUnRJefcv48uSS3BTzCIw7Nu0V8
RXv2/9VICiIVMFMaQVJexE+Ww58IVOw25uZ7jfSWAHsZRyyzLlWsLuTfYzseh1EG
f7MrIE3YEGxByy9BxUMA+WenVhAhMmbdRzBB/k5XP1Le9BRyww3GQEUF4Fjicz/Z
/Du06q+XEZ/om4LWaRvCXYTLOIzJaSJT4k8oJSGRQM+zjXyX3MeBnXLwLMgpiUnQ
JEXLVi1HuqocOdYur/2lTdJ1qpAtsst5MUMYpw2NRsSDza/+YgYVcZh/StT22gkJ
PpD6QlMi6N5e9yp8qj8T/FJHQvNkaR0CNtWOrJhhfAQNqGMyUYe/o9bB1OVlvIi5
2oYw0hSusLVsu9ZaYpKFSgy60G+PHO2bb53SzIAVj7IoEE81mREH7jH+Z8yt0Eam
z42pkLxeeM/ctvh5mBsLjvtHNifsN67ype3L6d8j5nYWZkKXI37kqCpd8zId0Sb6
FlTVrYhPt2eIepmL7N469iRQHufSe2WYQFejPwTNvq7TjoDgTVwgtje5SO8cGe8W
ES2VYLJNBcsxI4UseSpRd0l76zWoYr6S2fc3JjCaGAVTPSz+mHKQtlN2YCLqwlKo
HO5xw1RXgiAqiaTMiGJ5nbiYOw95HCnREPijcgLX/GspoiMYz59MREYUIpcnJN/p
F/6qjMLUXbx1sVwkY23NNRIQfUilFrn7/gNvZ3fo54ESTWbMm25lJ0TF2spI/GVA
NBO3b8OptC7lA0075gksuWsiP+Pt371YEzYPpRJO3+GGucnt8qb9Yr6uAVIBib5r
xT15lyBAnb+jGEOaoDe/xTalYN+Gbe3pHlAlT/veJqF69h6eoIwBvgoZPiUS3czm
kfxd6zko3fN2WwQT+DUJXVBpT/SyRJ8da1Cep3V8qORr8GuFmCUuoG1lGLxVujZO
bzHHjPz3dElaszz+Q3zRWJAP+yHcFAbbbkyMtUxYraZ4+VWzEIW4o/k04R56Crrv
FBPpbQPJ1m4XdWDfA9Q33B1D1bzTQMHi92qAx+AGDXGNRs7al3RHY9NgMEZGxGk/
2keIGutcqt9v8FogfcL8+JiAYz0z459u2qZrm6gwLKIOGFdlL4gCIdy4N0iAeSIq
r9E/Ly/U6jdPDeneivq/CcA696m/6FqumGcq8dlmywQ4rqY9FA9fa6yozEkcxJVk
niMh7O+N1lsxk7ZxgHkvey7aXYIiPVL8dFCIRBEn8lr+DbvKAkeTgASzScVQA2DB
h/ZT4p1tfnzRWHAz+VRO/QIcikUUw9DRCsbpQK6ojdMOojPrOjDiLj0UBqbJZWmB
73yUlhN63MHNKsIBNDEtRGZ9imoVjwkEBWr0VA3yEaaWOkSrIUrSQca3jiWGij3Q
pfZwYJnPFbiQ0YH9GuVCb/BpsCaR3RHA5Nmly/383i5Rl1RAnqbH7e4tsIPY4POf
79DbcYC8lOJvE/E1ZbCM1+3OFRlzakjmsw6w5prtqXP+rqa4mURXNeo1PWjHuCkr
SWEqvhQKGjLCmjmgIQGstLtU6jAM9bxTMZ3VUCH2FUr9LuGP0iIOATKSHzbcnsoG
u1tMvZlH/WxsGaJ3PKjqRL+y+/euZVy1yd66t7nHfKvgGF1n8TjN8F4g1XKx7IqB
2Rv9Ip7Hby+6RpcAMFWOp/ekfO6+e9qj40ixK5p9CgWJVjduXYvyksq9/guCQ5u9
TIulIFR4gTRivgnHji7a1sKyZb4YDbinONAnBdP9skR/VjRk2RaeIJRPdu7Jm9yU
LThdWb820od2j0YDZdScgTs9r0eI3g/QjKG4g1/Kz2kF6h4k+41l1T1QqZPaIEHP
WhIVtTHr6/28FuhDNp79Rw2XlE2w3iOV72zsR8zHnVfu/KLEf5UlObJ13UqSxSX1
gULwMNYVKr8zNkUqPKUjlzmrHjV2sLN3u2sewuCqKjucxW/aHmnkpeX0X6vQs7+1
0AQ2zfSFCG6JXZNPz7r+38TOb/Z/p9iO/WWh69WeP4mj+bJlDiTiKquaxKXSy0Q5
ZAumY6BNfIq+NvdqbduE+fR1xTpxtS01nq8eE8AVzbW4M0f4FRrO1ZmL2KjewrTn
UYfBuY+D36SfeoAtnPoTqE1SFPTq1yDFTfkd8LY28OGEz/BFOvHcyArXGWTJK+gy
0pEJQn1ZPpJxmUAi2U1juhLFx9kmXARGXCcfmTV5+W73txUuQBYNWyagTVE7iAdL
uwbQfW6c2GaJLneAWQzHaIrYJm2cUl1AluaQIJrkyxjm2+wQ2EQN4wWHJ6WhEafI
eRy70iTlj9+VcQbwFQqJJVkicBhih32Zr428k1IPzVzywT2vzAVFlLix8Il0WsUX
vKw3FC5cx+1/4fjr9df9DWPD1MFSacZ1vf9qjJIwzyKUkI+nXkbzYF+HKYB3QW4G
8JwGRzNku7NPJXLURJ+KVMyu99KQcw1WKGF30gsans0McgbpOMCsAeZTP9YoECny
/mNRg4/Nshq+nQfDi3uudnS9WaEc+csF9UK5oZCGKhYNuLNhfswomT1y1CrHk4DQ
KMB/tnrhu0eLIM68SZ7alAJ3U2etN26kOQMhshhaPla0n6POJ13PeyW1Z6kKszNP
PdBe9xv9lF3P8C2rj4CycfmH30o6eWu5An489FPd+0VcXmvOCL4y4Ms045YSQpqc
k/Hgi7R/IqNzKtzOl+RYtYZIo0JuhdAGJyrjC6DCK0YfTM14iu1/5ZiwrXniBI7d
TihiSxN/v6+01FBEj/iJYr3S36IpFZ0m4mIcYqnNaaR2SvSuOXPxemqa+Qry7n0l
Ces3EFKvIT+s6C5JXAWmyEq+I487sfu6GjD6Wh5saPQGCydomo7Qv6Gm4WF3mwGR
RVbVKmuVM3CKiz7YWiL/bk4bq0Sbw2Zvlk6vIC4ifKTM6SbUNL8lJDE4X7ULgsrM
YnfxucgIbwShxbGOfr6tAeB6qVy6ly3A/gS42d5BFvHdUmhZdn8AjyoY7ET4URaw
4J9Uutq2JEOp0kbiOLnCuc/GjkukhV0/yv1g9i51bVmIXjkJnl9ltZjGLcsZLNVA
TgdZhKq5ojA+I6Me+YMqsRczO2p+6m2NYe8EXQH4m2mH92BUstsAhfTKoe9Lhvcd
4LEaIsLWfucftsP1Sr9LTd9nYvSKKVRr98TxfYf/GrP3pMGQkdyaFcVeSqOn64tl
Xhb22f1hSYrkEz2eqampJRYyZEWTmxPRcvqrYJ8ta/5Sds2A/ZiU5E42x3nrZ2BA
Fh6+on5oavYGBjKNItVr9xX2IpU1IVXe66LXFcvz5XRkjz2xP4lNj7k2CAk8rRq3
apNUfMI30QE9odP64dRXmJh7VeC9Ez57AvTvoBaq/fkcLGctAL9dXXFoTX4mrDfe
3P4le5sQwU+cOWLX8UTlGp/vfRgtqVhDgX5DVbgLzsqFpijXHtnQki40M37HUV52
Xz1GRkHDLq0ZO6n3EDcdZinjf3nP9tQXphMUVERmmwBYb716c9ww2jKpuBs+a1mu
avuQg82pppuUUXQNI0tW5UDviOgk1BBN5w6t0ChrFmEK7Z7Yj2nbJJSJGYRL1DVX
giR3WxpxOVEmlEOI0cRVwWaz8XxAyyjvww+QO1FLZBzcuOzvVtW5StM51HFSwW8q
fMw71azJPzjnQzEVRLU7tpYDEEOhihiUMuxEEx+h4GIczU7DBplxfSYb6yibMshM
x3kX/XwpUziTaIjCc6c9YAOFHAwGX82ztLmA2zAxamHM5IROUOZQxSu1DN32mYms
RwxYxMCyFUDkTYYmgvtka8fBGGylkKbUQszBsWs5bAFY5wE7l0d4Xx0aynCSWdxU
hQba4JR0i0d8Ky99bgR0oaaQuC8Faj9ivz6q8e/F38eKDjuufxgZftICS9FeQ26y
sI9XCfmaQQ1B2MO+yXKYVNzM5WevzNSvgo2lO5oOHuzu7RhKOOqncYqhgvjpXlLU
wk/FbwpBjF5LwC3Qd1Lr6WNpZG825b9W/09STKlgiT50OE6wwg8XX/+l/00t8gZ7
Op2W2lscMMygZKS/+/ktr0KcaxSEI0HsE9dSKKojhj1FDeGieMJgEQ4/3n/Ie6lp
Mu+zK/pGNJN6QR+ThEjdnrlhvdCSiIYRzkC7RhLCFHzSN4QI3gU0nPIzF7zLs8eO
MP9BtrRzuEMyUXngKCOGh0wQEQBKztLYU47b7JRtSrtWXBOiWtkTVq3/e425Lsrf
3b8ZXH4FrarrbEnipIjpHx0ywXhtM1IE37LJSoo1pxpJlW9bpx54rBCBbhYGJCHp
pQBAmr2URYQhMR07hdxH1WD+v3S2eqAaXqqHTBi7+eUU8VGvFuKWC3N900cxioom
cDYXU0TEM7e/PkdFJ6hpFv9ebY7hQJPO/S4Zb/rkhKRwAtl+gm8w2vVqD05kf2Pv
SLhdMNoIzG5WXUXyKHyIXcyQ3q9zjHX1mckXJMLPflHzCOnXG1A8oTc93qLOFdiq
B1Q09y4J40m6NcjKvJKnZI2H2EFJs7jWVqox2xko39i90VnCYbm0kj6RyDXB2gUh
dANfnNOjZ985LbFLY1irYAmVL2YNnApmavkdNVqP24qI2Gf8/UZJPusupUSrHNgq
6tMoYosUaBaNgBC3gHiaosWcCFrd6r7sGWb5T81GlhHwHQodYthUircvu4R6L+LA
a+/76ByRKgITG0iIrCFVzlh7S3zuoG2jSL/jUjOPsxa2QAgUzpCJQdFDs66f2WKw
VMFJFkl/BykMH6RrY1AhCk4zaThUjJaIEMmuEP8oYsEwCvAld4ZEFVWIKxSFk1u6
QivvUq+AfL4aJbSO33j7pZBqFphE0FOhMzTxu/E1wM/dWpFVIlJZkNlVGos5MZ3l
+db4kX3OUsN7G8ybZHpdf+gw6EMkREfqcDLpzZbqbTNv9paR4R5qbw5HnLR5eYIM
gOrTCOGk3hhuhCoYpMKVcoGKs09/qDvm1IcOQ4HQmbdgWDPQhENuWhwf7adS/v2v
Awd3Ee4IKirw88YirSq/eoQIMV14HxGWgm1Glcxzcb+AYf29eVagtUBoGBo3mKZE
FyRa5MHaTvyKTZPr/KsptTDCmtEvt+TRZcFWCpIYn0ccvna4xe2Q7ndqTU+yU8pb
SlshDLfL0CqKRZl9x8tei/Ka7G/O+t+QzAZ9QoZqIhQrkDId7edzIX+qMEb8xJjs
ykYyTQpHsad81KGLk+AbEzHEq45nwiRgJo9Q7qIgxZjjKjMOBGGHNKlsyJu/k/BH
AJ2N0Em+dqKVQeJhdxsFutVyW2Y319ySDuCb8lqFYeMgX2vo19iriXzowTOhGkh5
Tv6d/wi77gqKQroGc55htl3J3YU+ogQqDWWgMHe0R7OIA1pDNKB/FA1lIVeDMk6y
eXQQL0g6543HpDOzp0GIW+R7IPMM20P2PTv+py+wj/mPthqoJue5FblFU54yXmlM
MO6pJyBCW8TRf5wv+j4p/4w2+BhLJZlRCYX0SQhoSDRKJXkUZJgoXWxwLAAdLXeU
7xOj0ayWfsb4n3DizC0qzoXleBZhKtMRmDapQ1RwLMihvOEkuul9Rz1TUaVgg7PU
L8CpK2krlIAtI8h2p/AB55p003/1ackhY2/uvMV0KyNaSRqr26u3fi6GXceQS6JG
0bjbT5BTewXbfsG2T8yl2H2uf4WezsMAUej0pMUbZCqOAsHutTX+1zqKs+hautRS
gfeGlns5joGdYefVrJxjg4y3jVsE79zpSbaybFaqOnbTG1u3Iu6xsuNnBQbGWaqL
LmROcd12ggCn81AznonW8SEik0FgT7vfBC99CeJQKaTXTU40uaQtomknO+17NNTf
au4Rf5HLRcmD/XBqfU+2aQogwSHmY7ModYGASdMGQLg4s6DUdrm1FLqQfwR0zNdU
QLmmXx7E2EfEtwDKncztHrPErPSHRxUEbOMpvOPnk4DpP0jYRXC/YKFKPlCRNxw4
7jSPVbVs/jaI9e1GjBB9S/VTBTuIKA+eUI1GvKhyqOe/ruoJTx6BiZV8Rgd9L+jT
XUyX/hQpEXI3kpBmFzwlobrE/jde4y/8yCYPmPri0T67HtxBJK6L7SlAfjn5Lv81
vvOLdlHTdBnCCjjcWkEkeW89qbXFVBvS/3fPakeZTQo1otq7NJxHU+nysGJVhc4n
JXXW9lIwImt5lt4q9inU7P3tvASJt+AT2kH87OAtBiSbAaOIxLUvgbdZ9t6RnZE8
UFtBj6J1SO7lXpi2wRXdbAwRbo3h8GqD5UHR/7QBR0ChPLVqq0HhQHTxktrz/7De
0JICQSDEMr2fbaEtmsIl+0feHMMiVuW8r4EFBrdsl+ZDsmvvayHtef+Ucm5ZNe/o
b7kldKuR8A+jkUB/l7t/sj10eO/r1qHXt9zS4VXiQRMFlus5VLTcMOVEqXEBfPe1
5cyfCMEH8FF2wxzLmTkGrrMC60H5jcGCjSX49SUEAMELT1HYHw6DmGedM5L/p6wz
orsuP7S7G/khSFToW0qZ0uSuCYPIV8DzB9cPyrweCTSbsSxCv4MttB62DRMot4xg
PJSCWCff5TkVBgO/IbOHcuGkc5FhhEqBr/bvHY16k1hLVJdIfrCe+9GkGTP12Bi8
6t7i5DIaaViXnBwSWht6vRERHMcsS/0uvb5hmpMqJRnsrQdnqy6+xg+S94IB7W2f
nwORDN5vrAveZzEpGVk0T6+sVXGLc6Cj3Kd89IspqAj1M84Vk8mQxynt5tXUYK4A
LpKi8Mxwm1VEw4EeX3M/XdOpc8HfKMwCZ94gDEgkOOxuSGV8F+asPCPCW5I13loJ
NvDIgyVi6hmSy+vBRSeIN1tUDR5AuHS25KNAGhS/5fq8eDah2VHcgrb3U8Oc1zvA
bIzb9lH9T+j/VRdnThnQzpywMaNcHmBbM12Ob4us6RiNg3Ms6G58vmfExFfn4QC9
i9ONSSJqfboWAEK5997jWYXnc0e9pJNMP/MgxfYsSvvxq2pqusmheRtLXvWRSt/q
/NXVHpHh6wIKVO5pPfyYu5wc1HSRD7tzmbF3/gah0vQ9ewUfsnw9AI/SQKqS3mRo
kqRtrBISvOXkYbbCfqL48itB5Fx+RCPJg6DxgAuGG3j8rvizfDfg1u/YxvH9rZKj
0501+EDup37S/jyJ8KKzMFIdqwtUFRhboS3dD21ANB01cpblSRzYNXf3B/WQ+XTW
XkGm+s3ZlNhnWu710LoMC7hrKJBr3WQuyFMwwhRM7FrPfb52yTwa9WEXdY9DJBP2
jfBMRWnSZlvShx+tlqX1LxTAhGhH685uFcsPtERh+8GYbwWOnNVxDyvf+K2g4TvE
w1bGZqQwXDP8ziaK2JaPcX7xevBHql7tBg9GDb8WboadGNdeNuwC87Dc5xUejDx5
4+/QrQpfzwzu+0ImzdudR+ufWhg4l4vnKcHbeYyyrM1LH9+02rx1zVnN6eN7Pgrk
OivksJ7RYYYGK2sYZ+tn4KLFmMnH4Cq6ohQAPzKIlPwYGJvxI/32nhf3GIB+xsxi
cTKtd7GEN7zVKp0JZQdLUlnL2+9YEYada5VYmASA5EEiEUNXXmMfWpFkb5l4Kqo5
3c1D1HdV0SpS/mGPEVwY0GUwTFP13ln5IhRp7coVxDMOhl1IS59ooAuLbxSYaYht
hMwD7zcqT1bpM8Mk73e+XwWZ1jiMUCSUUw0TyNxviHAqV56xJfcLIGHFOMC60Yk6
4LYLK4biByYCSdyQM0tP9yJKihhIAqCD4iTn1dIBYY85ursXPlNpg6zGmWrD8hKp
bp+ip4yUx4HjsUmVRYVXOs1phhHbIBNTxXCD1VwzBwahfjyRDMXZa1Nqa9QJWEC1
dgJndVgaEY1J99ANQ6DG0e024NuodO9PfsDKqIKuIa3awJP06UslqBA3Q9Vn8XfN
6pmxfUGmgF3cRWi7XUyEjrH5BalAnJYkq/lxsfHRHig/tgvFr6XwZL8jA2Zuw2UW
toQC+9vDL4Bn3UXFTvoqvsCKUUmryARNkCMVMYT0OQeJ4n50jPe6Dp8xkQsAQ4l3
U8BWM10pteyoAeeJkSbmQ7ZLdFL1L0/PrP1z6HOHY59lQxTaJjYr4arB7IZUiQiF
dXptKAg8q3jPZG5JHfPCKM445MJQ6XfiQzvh/OaUZEV0Bd62Xqu0iyFQpjngZjxH
Ipbn2j8RlDo6zBJL82vV6syj1/J+meJxKiYo1dVnabnLGZaeQrioBFtakoRU+rrf
XBRPq2JKoAKXr7oLweleVKXXzWe0i+WS49njFYmgyYjkR1t5XZg2x7C222msDpKf
LR1dmL75WyC9/sEFemxcvhOyM8k77QdeCXZViKTj+ABgz2G1/sck4YamDVbDiuBU
eBHQt/1z+0P0HBrRNYKsZnxZzfBUd1u5Bd1br+SgtzLHZh+y5inmndgTze+MtrrM
K7OaxZoTT9bLHHCJR3biCDDXVm6srJ+RwxUSER0saA14GERkyOJO5sGOKwKpf5Ss
PQ5smh6R3Msv/pQH+qnnJP0jCcntRJhD6Mp3y3RVr2WNHz3ZATAw5KAePH4Zht7u
7rLAJGdgRmUblVkuPo5CipCCxsVRkGjIr96hkqVHv3LDp+FjmbTUyFf9wQAXxbrM
w0w9sb0g+pQZgUZNa19MHeJwFhYH7Px22vj0BqyrqYbR6CfV31XRfJOuKII85G8C
sz1HdYcUeFmPWpJntlcSEdymiD9fw5xmOZ3oFVanVdd32VWbdRZJGjYzodkqIgRv
fiTszpcfSePeu/S6rWBgmFt4J6Mj3UPVSZnUwrs8za5dNKh4yP+e5qrWyFzrRZD4
Mu7DQVcb+djAD8s0NJ0OJqOGsbUzGoDtk255zN6KXrhJnuLinOsOuujk7Nc7cZ7/
Ios3d0duX3sKSKDassjzb93pmECqOBOvxIS8wi2VMLlrdBWdbDsSFshMQXk352qV
Q4azZsVPoQNM6qj+cogkVJ1Bz8u2Xur8SuH/iitIFpWhOi2ECEQBAvFh0FRXo6Ae
4d2D78ln4ogPrq2zI65ocQC7EG4TCuwmhGTM1EsnaWvcdqWGKtC8JvJyiMQSavJH
byM2UTsTiVPb4d1O+LZp23pOX0t/xIhYOoaerihrr32vUm/jCK0YMosVAuuw41Mg
s+ymIxOS9VQ7WLJbYrAJl86ygPNuKWJYR8u3yBBkb+gD8RXjAgfhbjQZ98MjvpAv
+4+5DDIKaZJO2K3lMFqdioHrJU95ddgkd3viwdui5vjrKh6zhLf1lT4NJfPxXw8i
GNEuVxkWY7drjKBzku11n0lZB0UPFyUtx9SsFvB6JuenFXwQiZEf2/g/pZqhp250
RtuTl/Gq97lAtbE5Wz6NlapXxnG1WMgchVpngGI1jj5MmVM+rONNwrGmuoutYpix
HZRoJP6I7wW1BRqnrvIf0/Q4DEWMwWyNjIJ7fsb6Q9HVJsShNCYg2/U4kA5RocEZ
kbK5Zg9KnVeef/9suIOdOW7w7KggG+13EmcJ/zNBaslpddjtKKyeEWk1nFmOAo3T
xLjdAD8ITbAMad99dYFsXoh8A6E+W5MLCEQy9/S9Ia7/Rw1pYyw2XNjyWFNhRP08
gU3T4pZ6KozaELB4VInU8z8F6FPBW9vjHQ/CliteyOIImXX9FvBkNlt6mVnRWOEr
jwGnC44aoxoJQSxtMUhXdSN0cr99zlX1+UldX60p8NrpHBSpSw7HZEqfMV6vEvxw
0ODxzIM++tou/x6TpyHxr1oQLvup4SM5OYdD+9HX3vxfppVnZAG1Rpwu3YtOH1ks
1oNzyRtjVPpGJa9uPX8S2Krk7DaXzNIcZSqUzFBYfI3DQPpJGovSNSmTZB/VjkMq
VbAoHEs5OmucVVs9HMngVzOWJIQ0vWkSrA8pmWejajuxY8BjUoAq+X2JLfZ8l4gA
xohd6DClb1OO9nqY7jFO5FJvj8FVKy2pV+XYxaqA9EiJpiOYNhoAYz9K8/OnyUKR
W7VgfINfi3qYrMFs2fu/6ZVcB3M0JzxEo4FyLpeeuGg6zMP83eP8dZddGepv7+XU
h/hQ37WMm9gqc50e3f3SEsnNzVE9FeD07gMjP5CWLtTPy2cvRdZrQtmMb9HyX4vD
GEbqTMmjLuX8mgLMLxa4HPgThvqFM8bsFv+fy/kxPCMvtK85ldI51dbh2nnuynxi
iNoZiANExQIFuI8mF08FXlsu/ztEeMtSyj1Nr66N0kY6z2rR5Kq8HZ6tv/vLnXFV
GaVfh2fYslONjIEjEORf5LOkDpFI46m7IA5eaZMvljBjtHYl6IcKxPVJBwa768Wk
+ley6rxeQw16FtourOPTBg4njiM+W2YD3OdAomK78fEWSRbFD2mRWLDrUvuTCcQ3
MUr0tXb8lNFTU6+CILr+IHnLH1EOTU5Tf+ionKSHWF2CcDvhdcubf9Qx7MkaTJ+y
6zP26UASvjmzxcSuKGFmO9Uvs92pNlE1U6I19pEAyyurty9OtNHu0FHL4R+geL36
c7qGfxv5/xquGbVkCIX35Eg4PUgl/k7J/sq4WmmBsWakOaAJmYRUmgfncuCsVGD6
oiri+bMpa8uDMf3iouub8FWLq15D+244aUjwVL0c3LpXcSB+WcRAa585688Jtk4l
K4OaZrTNZOLLnMLYjWdlIyHy1XaCG3H+jIIn1gGM4fAdBq0JnXj3Tcl0Kd7HcmLL
3aQKXeWVeq0mZKDQ+nIqLMCLTFhSp3XUYBarHE+QWo7CQ/0zJ/IJyt+D5vG2U2Nc
8NXm++va7vlr7pADzT8Y/nRlFs6IhjQ1A+5zWf+yE6w/ieNypPA482w1ZQJfHGy4
u8JcGvWUtkDjH5aKXD7bvU3apBvPkTYsaa+vOxgn7q3Qy9GN64u429Tb+h+X4205
dm9piMdyYeLEheKX3m66z03hX6Ily3fiWObiyGpo7aaHv0PgFBH3+lN7yJakTgs4
GQpOj2cSZ2L9i4THQlqF3ltFQXYuSlQWIGeslGynR1C/Gq09SGUx3ipD7q/R9cuL
7hwH5wdHsGcIq8Aw9SlKwN9otQGKWts6TbdNOVebiGTd9PHebdBkoaYCpr45cObW
f2eb89EQvDXVYwu3GpkDaKfND6fXk5yf9VfzaqqvGXPOTzDZQb0xyMQX+lnb7xMJ
e8eyTa/CSX1x0jhiyaDT/g8GPvV0srUbZ8pbvOPvEfnW3wQdn4gsLTfWOVnTmbFm
Lyv2UKjPojzhl3bthqcPcWlXqv1MaCjQXOXDJE1roL2P8ycVs3kuiyJ5+FfaguiF
ivM9Ht4vadf1fpZqtXKp7CT7NS3fjwYfXfCVyI3/s6VGi7uDwwbyk0DYGIdYIGF6
Raf3T7lPpE5zUl8JBb59+Xc8zFeRFjv0ic47fq8/i0oYb2ccF8LqxOg1qgj24xak
gV82Y9ws4ddZ444Au1Qd7BOhcuyJLCEawjar54UtbmRA7B+tY+qLErcfrtylWVWt
qg0R8/+l9tYjKejszpk7jqB9Km8CFUHynVJhU2xGzHIG6a3rAohNpHKrLxdfLvk0
wpPx23Vl9mFVz8HJNrmzrB8mt1qnQDHUtuMgxF+Lh3qQutPXQhpoeLpNZb//hFMl
G73QUosNIxIZsfhOVyqLyc0I+8Dtz9oxqFZEfTZmzdUx4m4Hvs0yZ4ujG0VDWAru
F4UBq4sCymtmRKzAPo7TWV0GsmkqpMU+HXb/W07bbPhZq7A6dEVMp1H955VyYcaW
V99Z0nOqppKfTDSB4jsqsaXMdCYyVBlWjawCDgt51ZT/0KtPQb6q9GLCwUvHWsi8
FjfETPa0ADQZsSDv7Vs4hl3i15tKH3O/eG5wxRdbnyCz/POKcNyUGEVXBZvwo1J3
lMAiziI/Ck1Es/tyIlHPDJ44pPMoF6qnHXT58/n8/nSTyiGhRNFMcVIaBK7Ajgv1
WKpuBOUGs9xPJxTaWX99wFJpSkie/G18//bDJXqERz3l/dghsotwjDHYn6GZ+f2v
JR7dZZK35i2g0sZejLUHR4giFcS2bxrLlUmy7qEP8WqQlI5IgkFaOWR6t7xqVajy
U5SGa/auk4U17UVYcHb/ElqISlTuzD6SC3qjtfR+cpKtzDDtRa0Zsws0qFldpAIp
zgJeUyGKL1kjNkPqq4hEYPWtl5nguJTAhotKHny7Ay8KjEGEJ7JmhwB203BPLl6u
DwAhzwaPvHIbEHxfB9zBNWzSXPy7agb/M6sAaTC9LeTaQnnRT/SJ81RaIDSg/KZm
0WY+323ydP8+8bmmGxeqxbpUanThmXuR/uWn2QpU6Z9shGj3LDyT8eO2NpdmgJGA
622AZf6aVUBU7XqEdGrCx5MMBBopt1aHv4LCtKwqIoddqbHwuAY/jr4dVVdaamG/
HqOMBsGEWJqAtZp+8o4KVcwSuih7whoXkMVoV8Q4rFsirnIbYx5u9YAa0N5Uqz+x
1S8fIGw/6fP8El6u29Dn3/+dnuN4BSl+cdKdMV11v4jCo4wivXvhqttgzdBtFfV+
FMrmbemSpBPGBdvjABeS1tZpMIpWy/2Fo3y8zsq4r9u6m7EMRHHZgacmEr/IxeGY
osfo5ebGSLRTGLB5VO09jTcMNTOJ0XvJej5skIw1IuvzvT+KhsLBIHC5udRdxMHe
tqQcHYA8P7R6/ZiBnNxEG3BY1jrN4vpTF1RE12K/f0aB2JWjc37zB/xJzlNS5fV7
8PyTO4gCqj09Rl7YYyvbwesj7GHRYaSpx8LAwpbggDoLx8dK6/CpA99Sbug/OpyN
d1LxaMjMxhSnMBVYPP9ngwDbek3YRvN4yGRKwebBvbNyV63hhBGzLCamu3BvHgbZ
jl0L1JjvKD/dQ4mVtX99zIMzqu8hoKk4p0qNDyrKRGQh5TR44ugTzAZ31vWpRJCe
wQSjWPtZM2IocSB+ufD32wglY5cVSUIE9FdMNLWL79FQegnJ45sF56FEA9LbKPTx
tzL9DYF1JACud0W5dUVzh0h+Itzm0XyTebw8yho9ap+52E7MGVGQDzJtIcMx+0y8
LmrM3FgDzH3TiS4MZ2N38s/UGbdgGN8M/o2nkXo2fXrkWGa7s0Hnwe8IeZw8eA9f
TXobjQ5Rm6Sb9K+mm1nDS40B8AMRyyG2HYsDqaE1KOSPxkwt5EduDyelSLdVxLqE
BT7kdUlW/DvpbF49ugYi3jQlpQhH9dS7SU5vwrKFXayjVEYaRciaE47KJ6tzyZCD
h2QzGyHk+qUSSpH6kCMc7AHJMgOveQJHvzgNHX2aWjI1Az/QJl8i9+PBmt5J90av
x1iJCdnzmKbOMtvJ39u97sBgfdvADjE4l19ohLRBXpsquVV4Vn93yxjvIHEe59wG
P7rSCeZ/rV2aAfC92LA/i8ZH3hdBed3sJIg6f9c0uUSU56zdvTP9k2uXXDojsGSP
uTdGiW+vogdNGFOCmbQd8lRBz7TD/S/ez6QUauSJx6G3D1Ba/uWTbMBZCEkdUE+a
+NXU9cYzH5fNADUZxzmjGZenLAp91j7K7N2W8QG9b+kDky+4qm8zrGvwYHY3Q5Te
sCbltq7YqsxceiXoNp/1jbN++wGkg/klhVzT05eV3TOxDVTwU6OHjDrZsQoh7g3t
LNqOBhtF32LC9XVz1Yj2uHDos8Zo3S3e9u+XCdDvoHmP6FOL5DLLjJrseYJfF3pV
9VgXGV8VsNuD+TkwlHIwvBF32+seX9WdLdufB5LfTABOg/v8tPsQU0hg53K+J37h
Q/PgMm8oCfgBOVyQrTSI/jRKfa7MeLTBCWRvpQSgDgjXvWXS3S+QmY8LdPRj3W/1
AFt1MxODNuo3mIn4/9vGlYKe2jnTcpx+BO/X4ewjP8vmqmXoz2L9OfGCHhVu7T3q
fqatUexx7IaDtW4vtsftXIJwE8lHsgZF8RO5Ac8M5rX3m+hJrEZqQDXF5sLWmRFY
+ULeJMsLC7n1RzAj33dbNx3zOmFRNrZ96myurr+wIojUm605lpZISQqfkry3IGS4
+0sNM7WX9e3UwQ2X6rw5IWdQZmqyBnlMfg12aNdgnbm6ZnQdZtQZWZxO8FD9C7wm
PLn2/6PY6xeY5bt6yxVPwDgXjfZyUa0fIPex3yo3ubl3ixUBWbyv/qPNQMheSU0M
Lg8+VmWkiCQX3tKvO7vYXFyu4/YmIKNaQ2ItCkZaY06sY6YW1IWZydtwKfrYQDAj
xPSfmClAFhq5wlG0p9IYHMlC0rmP+zPJt44z/CXlIc8DfdqlJBmIPbg7VTvkdIzD
Wcn4A7onKAu0Ko8JRfUEzq/0BObbJxTY0n0HFlmxRoAc2zuUqFQKVfAQnpWQbTpp
aGXeiYsiYbfmgoDEzGBXxCPE6/seE7GPT4Xya00kP73OmHvg4Y3SaDWZfBts5TdR
qYjLyvPNdQoN2kX9sq76Q4Ta8yxBrL3z0OjWeY8KVW0OE4oA8hxbloB5j75AbOWQ
2Pq1jqewqfrweY8Tm/X2mzuTlDliIdJ3K7nFltoRr0s+ZlDNsevfCK8kqEVk/Lso
fkSDC0oTsxKRZhpXOFEyNxr4FLnog8+A7WgC83Vk0OhncwOMUnRokMBlNxw4qZ0t
5A3Uy/PDfOmynMu5JJvFDYrT53Zp5ZqiIp5revfpcCFf9nLcapi3zPn4NahGJ2jX
D25V2S+CUXVzi34HotRPdUlQ2ypsc78y1kBqIuBMGOym0+qyLl9mXH7d5LcTwYpg
tzK9aUDuoyHwb8ZlozPoXYvGmZyu1Mmehj3DHQ4IAPzrTX4e53OZcB/ZLxM7TZnl
efvRL+HMrtQLo/BaCZzjiiXKqAj3WVKH6GKiVhe5VjL/oun2bzgYAio0lVfoRMzq
vdWfkg7PAP0MAmRWCg8B/X/BjikX6tJjBcieT0Xhj97Mv9Kzx4/I6QaczVc09+Ij
9jd7txlxbwrnWRHQ/So4+VC4uyTuSw2SkCP9k2U1YB7C5bqfrWzh72T01ME4XmYt
ZoiubnjT+YefhDXxZnjXC/WdrSAX87NfzIfZcwxB17oVnvZ0Ajd1P9CMMsYegnpS
HiQRByOvqHgX4Fgfu+NDWG+MCqjkFPnIlDEcrbhAxNX3LHBWfvjQEBE3nuS0VFx5
KWXi6VI8xDQOOteaGYRMMvG8Lf8PgurzIdVs9KJACW8g9j8R3HnrQsTfUZppJtq3
AjeY9abG/GzdniO0fH3w0BYV4aTOrR+s0qJhg/5fwzxsnfe8E7dZspXJJGhIq+CT
ya6GIYW+lqwP25lrNmqror0dtNQi5k9a5cesVYGfP+Oh7n+uz5J+bGv3h/OtVj0c
1CidHuLSNLR6kpNq1Y2A9i+vCj03oN9l/7QagQa6uqXgo6MBNc6tEL5irSqGfDPa
2QOWsowqSzCvr7pQ00IanLtzmx/cPHqC4IZvti4A7v/m4dbVZLBQNq/utIqFSTqg
FAYXR2O1TXAyQfeYWqX8EH1y2MW4cq9nzDW/tDDRbQD/852WxLo+96dOIFDSu2cP
4PtSzByB5t1dpLCsBIsY7e2eAGjSvt1kGpjUVndwNkr2g+Ie5zjla6FGRLqxYLrB
WBQC9fDKzrY3YFf4aSzgxRwLx2Ljacy3LfDL8JxfTLUnSckx1+JtP3msRXkY65m1
uTDhE7akpJSGufGsgCZmoWDhR9mMYr+o0XTMI26fRsqcWF96QzsJwmkKP7s9cs7N
`protect end_protected
