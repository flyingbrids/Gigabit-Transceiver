`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
OWZG4ApffilGSrWKZ1DU8LRvrrHS3PeGUVVx68o5JpN7QusvCmT1mBfxNSt/TwFR
Tve4sVoPeZwQrMyS0ImdFOd3j30nvEWAtdRaV6mDPYHTABuURPyNP/Kuna8VYP9V
Ot9cO84jDhIMAK6xoDsnlM4QeS9R4pBPF1STeqKAV9IRLJ6cnRLLa1vBu3y+cgi2
vt57D24kGcvtM7BrkviIDfcITYV1Uzgk7prFKijnrZhzJ3XQbB4qmjThm42jkKRC
jLd6llH2B8+lucr5XCYwI4+gbVDnf8HznY4JyJgVY0gN3AsbAMGldchO8Tbq6L19
+hMzt1zzbxpkujG/1yHtmQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
HYU7ulVAplyNCSdwkPcyYIt5j0pQC7TGNjKrPe0OS2MlC/C2iLt/uxUoQMbfg2Wi
krW3lwdmGxUrVOuPwMP8kusz0JBM/kpyTwz+ihhDayIjLJbGWt/4IL8/tz7EDWap
f1jaLTqA/MhD+ZwTsJKQgzb5pMybMHdvgWT0uysY0jQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 119840 )
`protect data_block
SBtUvvGlrsnvl308n3GVBOuTE1SJdWTPAyqdBbvo2ADUvQZ3FvUa7zfPDtWbP8aM
t0ElYIKvFbRgTye5B3gPPvnxNoQpnC+jPUpleWUZYhhx77wb5SqYM1qoc9bI67yW
ZaLzhjT9NimprS2F89+BAcAAC0MrTZy8uQIoI0H7kibwQeB8a8Pc7UClMtzrU0lI
O0wSc9a9Reh+jMwebpdqd5rE6Csdr8uNkGnQIGZj42d/g04xgIrmTD341Lx/t66l
ADiaqsEkQ1nc9Dfs8/uSbuUrgti0hPJ/i71kqzSKgUuXWN49puX5mnxlaTvGsm5W
Odlntv7REAg+EHsiZYaJrgofhAR5kuLwwUM4oPl18d2c3LfVVQDOgCN4ATJE08nX
W/YRVWpp+UlvK6iWHUxIpJ+3CVtbwE3KQRYDQJMg/1loOdwHu3p34dOl90hBPq9V
bU3+6Kne9NWim0/xqJHZsbHu5a4Yh990F5YOk4Ftw6ipDKS+60grQXR+EbF6GJZ/
DTHfQVGUOg/vYSmHLSIZP+BMIgKqRu5lpehBN2p7AUMdMf1xCwDqkcgFn1+qLS+O
qKsV9FKBfzJCUlW0pdGXMn1c9+RbWWJR4TWoAKHR4kZ8g2ny0J9iaCZKpQ4YypSM
W9IG1z75GG5uGX/yvyYvJTOMH/q6TLcQsj0pcKmIYf+ZkL9htaRxs9IWTakWG8lX
AbHktlJTu8LGS3NY7yslNE2sABS7Xeb5gA3BiBFieP6OZoeFWMBejrh9C7klB4co
rQd2ig9KttO5/0HXaoihFnqYUSxZFzAFcO4wWbcZ5vdwdoptrvQMJ7Uty1hoJsWp
oPEJppBEjJziCR2U2PPTVLbfQYcYGWNxLKOOr+WsYm4qZeVE2pGGbS2ZyVYwzzmk
YxYq2RaeVJXertiZ4U1zZD9Eg3QVyiTDuxMBpnY+wxHoN9Z+cqz96BDMBl7Z8e2c
RK7/Ldw8lFcE6SM0r8z6wwg1u051le+fikQwcHzgCp96vMrZ7FxaNtJ5SI9OIfW+
W2ZKvawZYdl67GpEf5BmGGb16M/sT5xrU8Aq2+6suRSdhgMHl25mfwivGjAeV3mN
gz4HI9dRhLoKTYfT+JVAHDc6WleOuCRijHLe4rVm4pMLuNs6PxpNmW4cV2dWtaTY
5MUaOGWP4lcjNsf8DvFCTQ086a0HnD1XGe4W5wiD2M8XyuFsE/4xilBIio+sGGmT
R7Xun1hBlTAm0vALIIPrQnK51Avhvfly3r6++UsWJ17kjBbAND0M+fuyLs0Fl+eI
1pz6BX7ZjZgv68XL+F0f1mBerqsD7Km4bKxD2OCDU0yIjki3mYuD0nDxB3W20akL
kWakJdItXEk48YYK04H0Tg0MiZig7ewyD7usLEPmvf/iFXGvrfNXCnxi6Ok4R5Zd
gPtPTlJh/+OaxLlvhUzsAESpZXRzJVIyiitIeGdC58yy6/u7c/Rw2fcRxcv3dYrn
CAxH17kRyeBpY7CQl51am8p9V5aWhoib8Dbto0RXsvjR4VSEtx/XxI7AQkG/ztt0
2idiNwGDoxCh2/klB8aibNL1hLwEnISdyfWpNZ5G4d0Hq3fUPsqTm1CEBfm8VS+M
Okjm7GzEFhXKLYBphN8Eh8pAyA976wVtEx+iI9Jw3M56CoAMS+Gl3Pwr8mwDzw/1
8U1fHghVXbQKWdZtEyQTlBeEaDBA6L5lpU1bCscQUFqhHX3Ypkd32OtQ6N9CJ6p1
MiMuROYhqKe6xEobmT/MfjyrbFhOorp7qQNacAZSM0ZyzuVWOx9F4wN8t/0Q4xJx
rBScJqV/TABpssJbSEXhs7CiHXQBgXUz8n/X8gzc+FQmYDJSH+XY1gKX6OMwTG5D
4RY+SshxE7wapPYq9IhRJFUZiqFhsLLuzn5rrL/wueTXapyRoOodKfzKQVK+IeGO
p1vI9rpHwC08EBZ0tfy2J2xvJZHbtvP3qDdaiIliwmtPmQsMgQLHjL2aq9BgqWHC
sRicY/EGkh37oqgiqF0Q4pDAeIiu2pEVkma6Dfcjy3JjoIC+NqpxPYim63TICE3Z
DyvkMweLH1yuXxb12ZmVboJyMbgZhTC6rhJEYT3nVgfTszgoziA8VIZffbHYmN/n
3XNTF/tj3C6uCK5cpAEXg7yi392QtRGi6gts2/7OXOi5HxCUwdvZhcWKnW55gMlO
b/TEgFIuzsnvG8tfHB9IdEW6/epA/nUGv/2nIsduhnsvtVC7+SsY1sFwzH7AlWax
XHkMihuaas6ILiLPSDyKvg4wuqzz0IEUTwUM4IfL3f07WEZs/ewPL1CCHtA9rshl
Yi77y7fc9b+TdU+MXem8DV7yxCYVhpRgg81pML3vfbfZshG8W8MNYfyl/tOhKi8V
8wmPUtVzNW+eOipAU6VJNd7ntFICVHS1EpmiilVTZeUaN2JKMKH01Fi0ZdnEWHR6
P06d+rMDbSYiZtENT+XG8l/l0n7zIKnLnh8+CWVfTNMP1NWrUIhs2wqw5t0k3Cq7
hmwBfJ/BCW6YcjC2SHnjhC/uxrcD4m0p9HKXlahT8Iem5jQs2Yh5eNGySfUls30X
ILlj7GKMhPrrxYlIrfFpAkYDZ8g/+a3nw7vagN6e6jSWYHIFCkehIzbhutgd4tch
ilhjz25AuY+oyD6h3kTprbrqtqXm8MrRwvmXy1TlbIz6uoRP91j6DR2740Gc+YjB
4BygfWNfHLZvIrjH/U10ZqZ9VclIgV3ZZk7uKN60PogKiDzC2+iya470NiVVSpBC
bxMzdOA1Y+1DF6lGtI2FVbA0JiHP5vEQ96EZCZaF6//T9+EN32fPF5F4RkVzJzlz
U2dNiqCdfSZ7p9oA5HZe+FSdItgNkPecM+Ig5cl62iI8dkqvcRdprzKDi4La5+0B
drQ2yeZN2echUQ10oYNCiB4pv746RsyHPNbaMsNIkF+UoOeefEqkHSeJedqSI6LZ
graGMJsFqoMwnxJxeFNqWgGvDvvRTj6QcdHMGQSd92BbHjeAqlwZAQiy5/xgFuwS
/tMsVR7blwDnGSNLhmTqin+ZAnFpnLpQLVmvDhE/4TOxOx6h5yvgUC/wTjTCu4a4
JyDjxukMU1Kh2GWZgNJVoX51wNg4HlrAl14bxBzFUezZFTldBs767fhExOFZBFaQ
PvHKTFrt7WIejwhozfaJouzjgWZ04hu499sM4IGXeAMDXJNXsnKiyVwFOaLcrpTS
fFUUwIlH8sjAk5lnMkRvpha5hyxg7pfhfce47Mpucxl7YTiUgZULu0+HDiboyulZ
f0p0aInvdRhJ15u0skMSBBLb/iO3nqjgiytFwMkppfq26r4Hym+j/Ta5NLxFPPDH
WLDsTIE7ZhnI89USZR/Skj3uo9s688dnWgiSwupHoOc6Gpl8RFAqjH6FgKCxWFFV
1XA8O9aYHqgXfgHxN9NPKlHtG8dXfw17BJEiO4ZMKgukJ7F6JtZl7oze54o4jVXe
zUdRKA2RSygG58gXWxgl1QFHiMthBasKJ4L/qCZVlsxB+EvDMSSDCegDsEVUD0Zp
cWXghiqpjLVotvahmVshU1Z2V6DuJw+hlXagu42evO+HOLmauTFvTllpCVPLtbf2
BPHZhbaSCUUix1C5jWtrEdcDju3jg0uYuCf5OfwnjNWboPe8ki2wpZRU+wYwPRWw
2GPIkePJ78XVENAHhUBYshXWCBV9encZm01vBA6A4htt286/v8FaxskXU1/GV8cU
qLdfd7PN98Skh+9NdX6/KDk2Y8Jx13Ho2GE3A6c9jXgkGnlzuV4jKfJaLnaDMNhe
dg0icsLkxZnsZZc52wHBDZmvSe0HG6EadXAinmDAJed2uH6bR8cKYqEHGgMbvzCC
7OIqATuQmHD0WKqvWfyoFsmvoMHU3Wl6BVobg48hfD8X8jNbgk/LIWZ6P2Gnx7w/
XDyMvjk9mfbGeICPLII9Yk9G+WJUVso3iIusBEuNRVBk60pwrXYAE7JQx2bsFBwy
SxTiDO4RJVYw24kvYLoeipEAZmp0lB/qKPYkZpy88803HTr7Fx6kSXJXedeaRf6z
erF/x9bmDhcpKSQ6o9cP8oJlTRAHseKEpe7/b2aSuaoeG7TQ2Z/sQth+zvt1myTJ
5rgPYvWj/PG8C+UhhIb5wDWCzXflUyKZrUXns3bmYSpTj0u58CiDuF1vxZrfRwPi
Abt/VqXe5l2mEOTv+Kfooqk7xo0y4PQwaUqb6vjLElCppPSOlRLcj6ZQR6WfGwFm
QTOg/7Q6y+GxAKSJ/9QeGFRizYTe/CT5BB3AXt+uJOR1xSoy3BM8pkj6bqK7y4Cg
IxE5H6OHwTR57EdnnhoQ6P17dhQD1l5c9FxVsO7zCrHN14SARuDVJtL9CWF5K+qJ
o+R9/HUjGhQ4TdvRKfGpeTvODX2jUyAtQ9tYACO5X8Tl/4bBWEkQrhDloyJ2Ghgo
Rk5YGxzGuaLJuhPFSUBXoLMWDBZfuHaNDRvJrtdMqh3cKnnNVU1z+fd7rxOE9Dvd
HkxfmtNDTdn087kt3EF+SSF3R1n/vIqxDk4EFQieiDVgC3wwgLsaHs5kakJ0sQHi
/hNTzXBaQ2IfsGv6BpNfLnO29FdpVTh3wnarcEOivmtRuMpwv5z+sxUIUItiBvrx
tsFa25+nn1wAsahCurShboldNVQgwGiLJGSNAVTCy/nMqc9Q+WCrK6SOB4RTZNJS
X5A6wdy10S+QacFrSYS7Btqyg7/ngwEmMFJBIt4Lt6wlgFMZyKfno/dTt1RqUMBL
zAxBHlD7u/JjBZ58iwRofT+ZfBrMDT06SyBtKI0S3ys0FTwvch5zcX1uXo0wPfd7
lJXTNaHBodUaDKN57d5UcBqsJy3/Mfz34NsWoTie9xCNawjhli61zYshvvI+aDqW
QgXdIZvs/Uq/YI5dJElxNOsTxK/XHdIMrN8iO0srya6/aY3fDK7DK39BLi/Ivp1B
bcMVLoB0oRMmAsVlxY1IpmaG+IDMDncEu7CEP64/RkmQWeFDqeaZGaHGKdJ7Kbc9
r7QG3qttRbQzJhXoiD5RnPUgJbO5lw6Ue3JIGmB6cejnapv3SvguHdMLzqQmTZHN
7GWleo/9+6QOML2xrIcnSOlwGzBQI0eSJfE8JKroVt+bzPDj9qVf2RUH7ugrE4gz
EtDSfa472QNSk7lcLYbExzeZ5K93HjHwk0Wh/3L727I6LqXpgsXfEy18AIAuvteC
3rDKffQ+r/ncxl+m1yMf9q0nxQl0RqJ18fSSV0HCy0X1EWengHpWkN9gy6N1N1l3
uFrBrCWs0I49jKvP4jFjTgpTnbzI19q4DlhDbHPYifNJAwUDyFqTarmg9250SlF0
v3CqnVSXhvHtGf619tdglCasSaacUlv3lf6CxhCQy7LyWL4kSUN0UiCmDqgB074v
PwzFnerGIkJoRfA2RHjiChFpNw7TnYYr8ry7XYo/eF3EAzVUjHZtrgsaDHKN23Ag
7XxKyOycNYDoKk94TYmI3rPtpLyH2tHrcZny/R42/VtPp19+9E7dY46O1WCaHDZn
Dg8hHgGadA9UDtjVgmRxd41sqB56O6ImL2I6+8NgXFCI29X4jtFK09vMiLgozaHH
74IpqKWa5gd20DgXYYFEBHw8B8D5+MM9JtT0HfmsnSGd6ABVpdnQn3JyjfAHbr1V
zAnUNtMrZ46dHLYkC9sQJpf1favJ0UEDUcHfL7oADkK/FNtr0uE943f0kAdA2QdX
EfCNORIuy/44fALWQBIsPK2npku6UdPM8FL04KaeW1iMMwB7ly9qRKiVMNahbo22
CYehm7xP2kzRxnjT4Qmu/GLBYVjQcrzbhgVdGEqvVSTLRnzIbOKqbxohVnCdJXS/
WkGBtAeB6cRvPUK59HShLFV+tw6ku5XHr82e2rTzdb5Hc20EOjTG0qiMjzfm3SbX
IC9+npkrxnKET+caSBBKJD4+qaGOF1QSi7ZB/EhwWwo0LlpuJ0Sw1aU3dGwspKls
8GU6RdnA5JeEKo/tMhVCHk/1ixa+sasN+g6htiGiTDrK1ceLY7C7iaICfAK5WEUq
rZt8b2qiJJZdiKEXw92EOFP3NMjpcitAE4ykEAJzqMXWBblhJe74ge3An4csN0sU
yMjrfD2QCeP+ciixB3K8+g419VoDh3fUQoUo7EfiIKxzm/YizwHKDElHf4o9UW0n
Nl3tEwHtqcvZovYmBxFz39v6pJS5fUX7NOVGe9c2DZoMFTpFxhUISnlnbKsC3D7Z
7KnhvUfVM0YCrMv3+iKGo1OoO9Hb32Lm5Tefb3U4F2DMpngxF/Rm4koQ8gSRa7+F
v3Tli4OBBvmoqreYpYo7pVFygLWHdi420a6yjedkVK6eGfrpL+9dPra/+0ryw17P
sSa+Yo38d88s6f6aalbWwYECbrzaN+7oOeBiaiXw4RJL1HyDJ+ni4G+8x711aEf9
6emZu/QHbJyB4+zVE+XsBy1S5LB4grRJ4rkzRMfJdwKw1tnyQaCxwNJgAaiiFOmH
l+V4sNQGsMCoD+z00R5EnzlE45i2L4pQOrpon2D22fG80+5CYTB3KKX8RAxI4Bmi
pjd0awbhMRKguRh3sgNmjhhYKwFGDLxCuNaN4VHo9mcuQsMLZN1SHoi1eMS0H9EJ
IB6GMSnovx2W2/HhDtb04e4bCsekZfi2y1T9/bxLCM3KIwvWPEJrETXaS9S+ZJBE
GbGpyMJv3QV6faNssQCC7Z3GUydMS/lK4Tvt8kGL70m6wo04R/moJZKZRizmv8mz
YFT+imfrYEHi+JjkoOoqpJsYd3TkAmehVbt2czBr6pl1kZXUp2xNSpOLq610ayG5
jvNODpsPECfXlsjF9FgKtQYvlliRXemeA0fqp4zCbMb1rtwMSqcXjU70YrqpCiqK
0KExZmdOZco15/xgSwBc+jR8+AiN5o3S6pz2WrIwFG6Z43l3zpEk0C8Nf/uIYMvc
8fLJxnNJ+Ny6TLkzU+acqVAD0knkk6j9Z3A9CjnA4pR/tdjNl06pOvZpjP1qJSAM
WS5fbU0uVufmbynv2g6g3448EXKlg4YMIvd3bOIi8MF+JnDqHwo/TERIrm1i7PgV
UWkdEnnFwroFs3Vi9ZjchHuH/QkC47/RqbptPRRVG2PqenStQFdXDHd4jMoJNCeH
xetMiDwRmafu90hKz+s8xpnJVq5YPTI2FcxS17cMGxOIBoW5MbaYpEgoBdBA0mdW
/mE/j0IdLUO5V7VHr8Q4JpasfkcJAXMlBzX7H9loArfX2E8o92lyRXJJUKJThM4d
gSSaO3OcqmqW+7qhVSspqiocngFTIT8h66NjaW+aVfWQf/H8bz1idAz1qITZU2O/
qpOQvQNvjZX+GzzEmqhEGZ4Pjb9FESwlqMcA91xPJGNFqHcg6AjAYv4NqfB0rgEy
TV5CYWBJf6QhwnRVoxYO4Ezglv/HcdhSRSbxICLhyCRFd2gWAJ8JWbkb67wpn6aM
4OBt7U44y+iUEM1j3uFWg5Z5/ZH4PxS/psFuX2T4Ju3DY01A/UFGQQkPgKyGdcjW
EDseTCMLn74Ur2GINaBipqZ5cNeCGzxlhTlO4GNj4O4vl3WKGk3j8ZIxwO0LlM9o
NWN3OGkIiffyWqzjhs7ZE6PCAIV3UUxX8yElDh6GXqtpCd8OsKLsJPxlbaza73Hs
pg5QOtuOk0p0ncZPWUPEUXJROVDCdXAe2R+sJtZG6YQSlE4dNHn6H20bmK4vvjHH
hse5CdBYvyZFXtS0jUF3CNHPnUedybwrHmySXOcuXIV7+85VVp23b0Rn4WrETDjI
U3Ik6Ecc/pu3LTAtd7oDF+Lb5rAD+LkYlQH2g3sIhMlCESLJRSoU6oS/rXh2H2KM
3NvuOw1YoaxJQWiJnXrdj24cOHB0TqRKTwYmT9An9OImsZA6fS+EfyemzS0nndOZ
yKFXt6ZYuTSjhZm2ZdZVRv+2i3wnIWJOvI1bCQuhs8P39Gxrf56veR38L7G1jzm0
n8lnn7livG06k8TygL6R9vk+hC2GSUOnbEbNZLJqRHgikvFV0tURGDdqSDRyEPTT
XI44vZwSe3qOOM6Fq7F2n39MQE5L36UptRV5UzfO8Gr2/sU/1ORkyMsEis6GHeCM
REdinItzSkFb8nasnEFKrX3U2Zi2NK1hDpaxd6iDyzlpSuUVARMDJlVE1flzUlZr
mP55KWuEIi1316+ZsvuJzIivH7Zo6E/AFjadpnO2MmC57PYlebAqc5vHFWYvylWu
fw35+q1k+rg6DECWG2lghCmVhmslx7tKYASVtOEDJyIkg+8vGUQhoOkhunou2W2m
H4bvYH1DOUIwJxShyT8dpo2Af3bM5v8izY5HixXcBTekY/Qfu16M+mfiz1Z1P/kA
nZKFqGG5vRZLuuC+mTCRh8sumHRdgB2lBcBvLzq5h6YQUFwqBdCBYRSB748dqs5D
01eFHJxts89zfuBicbiFxznYRq5BQZ6DbNDf7gAnRfGN4Bnb2mMa3ck961UdmuwL
RDv/1F5JN74GDG0HAtnqvFbagFKfJlMgQv1alpnfXS/ub3UBFUpaG1JmpXFp2Kmj
vVMLodgeonb7FArqx/kmKdT9OKaaYHNaXbHNjLqAS1e+WltVG8ESjn51L3ZI2Lo+
uGmJ6ZASfBRqK3xInwokbwalWIN6VWsfD9EvtfX/dKlFpgXUu+oNcIxywzYnTlnf
hD4prwO9QP+xsO9fXTTn1SED/3/7pZmvd4KE+gj8wN+ToXHCKi434x7kjM1G9q/4
9J1o5c5DV9q5Sb6yONcK5kIkVD6tTieQIIb3XPsnYT+wl/D9tnVQs/IHmN55Qttk
iVqs+eBUyWcq156Ka71CEKLW5odBVQQHGHjjE/b4YMDGmNvQrQmwr8AhEObSbtjR
6zAD8Xz1BNyF0+dsMO9JHiRHHHSP0x0OTUfPcvc5YDbI4qjsQ1GaUKEV5JSCj3Yk
yQTDrVi/Birewk3057YPbJTecxkKioMHqsCcJnYhSxdW2XX5TNlU+cqxgsTIh2EU
2BMy4SAX7ig2tbs8Nf6PKg7g4tMMjAHMReB0b1T5L/Wc4d34VzU4eCX218W1/7Ll
wzApGXSSYHLRu1bQTdLL+ZP/az0PEQ9C2hgcXvosH8YlNtejBQ8RT70jth+j52lK
8wY0gPj8o9HUwpXuqkZPDVwsC23bGHZn8qW40OQW4NKIgTi2fzKNFgjjnUP1jRHk
hlRw7R1kL7ULrvUMajVb70w+ci1dTkHfQQ+qUg+FXJsoDqLJ65VXnJCtLAYH+YPs
GOA9znP1ngQYVQTFELEmsbZHXruREB/+gLG6Rmc5TSfnY+t9MTbQSEz9V74zUtFv
fQOFg/HxVbaNSpjNbv94YND3pw94wbEMX3Dx8aF8dL2OoKycMNNrg7Uc2T/gsuij
A7WV31SVRrQ9HH3zTyugbByf0xyjYCwOmSbByKfBrMwljKMuiDj0CW//HAsFCSyX
krI2B5zZ5w6heajTrrNoO7uJ7sfADtxlktO3S/1UViM0XeuQwIeQSU9lK/h6hdK3
oFI8qRD/ZCNN4cF8jCREYgNaX2hVwMhVaDtqQr9GdfHj6QuIdIEGj0oIDdNNblCN
LgLaKF1tjB7hzu25dzhv4Vens3jQQ64EBlgIF2H7PvpQsWreroHoliyHY8Oco+hr
eMX7BJwnG+dfRmxVsUBFfw6Ak1JZECowOYyWHdMRp+KNYgMofdxsgzs9S4hSe8My
NyphJ5sN6jNdJKLF7YXdsdz2yWNW5u545LR/MtvltHzt9rlDgv79zkWWjbNsnciQ
l5hhIADax7MMY7ZryRD8gQbPlokxm+PW/vueii9KBVTtfbtHl2rOzkVWFcozORf5
L04nIITOUUSFrQG8ZyvuKEEmSCqCi+5pet3lH+RzH5r+qhjV88ZF1fg44PHi8/Wo
BwuTAVtkAhC4ajGapAVLlXzB9BtFNJugje2rW+Oo72N4xsZ/fDEvMxnDrKNWo+xT
1HK8sL7YCTNrHOrqYY6synEFeERtNNQ8TAeviDUPN2SmwACHEZi+0QIGey7+uDVU
mVNDc5e9hWQbpmr2dwx+3MRsBwH+x3H5D7ps7YFQ/fGUs5solU/B8x2H1xq98L5V
zLGzbdQJavFwxHIqRTo21LAs0lKEx/B0KYgBewQ2QSsTfyMyL6i97bqH9nBkpVm0
d7HWmvbQsaOdiYunaSdDRMtr3SpVMKz1wBvhzXeFbyLde9a3fqTJxhIBHZxhJZDI
epN9NXQecw5y/UHvKm+lud3DCCEC+bIB0R8x55DofhahVf1xUjSSMSlc+bbxO6qC
YHrkhBeOBRLdrif21YwDF5TXVFJvfhwZEBmE6jsZ02NuKHO5bb2YUDCNEL/m2VZv
y8Xe8PbaueiU7WjGs6qNjwpg6HPb1DvxN2+VinzSCugg6TY/9wdSVCDlkjjiaUzD
cSCmep1uhH+sukFVy0twxT50gZxgzUdruUzDQATTZq7QJPydPyd835qd4hlMAq9q
+7+V6NEQw3j6Mpoj04x40xtBm+jQo79o8g4LIcekrGS6hP9WBA7RkOWi0NjFe0s+
wO7yZXEOkI//XrqsUZ6twtSY6StZEvZ1IA9e7yjxFce2t8ym4rRarj8mpp5R3c3f
olUDzkOADuRVTe9iN/F/f9+S8mGtCrXxXImBy2I0kOi7+yLVftpHIPddPKqPhll5
xAcGPYJwrQohEiX1jBK4Vk2Pcrz6t1HoOD3RPtlJlFt0aG0U63Bf+Guj4WNdIpYe
+nW6fu0RftmyKjhYSHZtlty24pRrasNh4lsD+Q+vQRAGEwfc5Er6rf9uMw4XdG/Q
TOIzojAYwH9+N7jPeQrdG7PgLAfpD3aswpVTPD0r6DIj/d+sypqrb72iENtQysp1
X6iBTeqFDm73ocjYvqk7FB+QE4Z2HgEXj6jp2FzwgemZSYGaA2FHmOKIFjjBMPWL
Bc4MEzzNCtTSIcnSZ1cvviQiMDzgAh4nXu7tyIOsv+SdTq8fiuaJ9dymyEuuVB1A
ZNXpsXNpv5CVU6f6sDO6WoOkJ36NwU+VC15hcj3FAjSazfOw3MlYe0BaTKVkdhhK
FK1ZSQgKhHo9cuBBsNu89Hg6sDEiTh2yrolMnsxVu5URJmRf3RTXQ0Y4brwtV+3e
mb+alhGzU+zuxpJO+ElLGGDGC/YvFY1L+OqIw+z790Vs+5jg2dMPo83itClM7PCa
h7ZFybtGg6hYjOCeZGDK6t7Cxa+KEqWmJrTBCQkuCQCPg+6OTR0yIC0HUsBbjIss
/8YhBHEdugKY9mQjlnx2VM2lif8VvlApHPrFfYjM/sHEculho64VVC3OPNaQsuU6
IyLW+X9TRXu04RTWgWAwMldb831VfGmY0gL3jSc8BHz6hrTH3m+CnJ9keAsHe6Bg
ti74lxGr3N2fzQc75Bee2nLUDSX0DxKP3p6+VTJ7D8ppR32IjXS7WWVld5zU7FZb
yhsx3yx6/nqKbe7wIbv9wDqAt7njdHqBOFsB/1YvCwoNSRkygVY5OSBg6SyCIGa/
93otvFtaNA4qteDEETEPH5OqgcrYGIuQa0jM6eHV68WztJrgZyOXfbP8OjN7qvn1
otrQpPIDHau6/YBXn6sLUeAkxANlQYC2LdLb5jWQ8ZBCaNxJb7H7xuNcKbLfYq3O
VGdwulBhjI5J5Cnwtpd7rVi26K8eUOdQXnxewmiQNOlL46PyNJm9Y6XMBgDNsJO+
6A2UrU7fpAS1KP7GCafK8thUF9ptJr/2s90zbewVO5u8o2RSfyVuDJUb5NhlvSBa
9AmAy0dHtVetteLk6rPvcNWVJvkUzUXDwy4ZtH/2BeD9fqa5Lzhcxr3G1278Iwc/
/V/MgNFr64NOBC69pt/4QXFZtiDaP5QauFrVLpeRX8FMbYd3P/G/8okgk01hAvNj
Of1fZLmyghHAR0lUWBUzXRKMspN/yVEWMTNWZtzMCgBDZwWFmZ7IeLMHkuvm5sd0
oJZIN4vtqNgAiw7sYxnDlaN6cdrY8YhYWgUNDp6TJPLKUG6CETr+qOnmLKzOXvB7
eM0zxA/wV4HNEzRP7v9tNS9TvZZGfQ8WoVkqs1AOUkyagyyM4uAw0DJVBpTtEd1S
1C6n0lUY7j7b98NBOasLYWOWmyUTNW/ffsxklJX75Pr/WAm0PPLiYFi2E/1vAkJy
0Jl2cz4ZjEk8Jf+2LAZYmdjj8nrhTQ2q+WoPpz2f7b7TRpvFShSURsAqXixRX5Yc
RX7IguISb2InI6+njUSMS7pLUUJOjRZ3T80yNqp4Jx7bJhMN+TZoFC26yCyuoxIZ
otHLm7XvdyDipLqYoLxMfDT7AtoEG99zYCtk+ARFAPFC2SlU7MXch4Ts7CogJZQA
VxTXdNe55APfKf4HwRDt+D7Vj0HFdDV2EYfpqBGHKQoY/DY0tiV3/Ljq9dAGxkn6
azy0IlEwh0gq9MX7S93tYg8R+IyRLW4WxWBhmJDd8Yq40WevBXSUquQ0n0gNUDl9
WFoVp25WBUNkFf8wecRCoBmmaMMA9fivHfxggjVRAgF8vD+nZuepSDQFvCx0zPze
rulwffNL6lKTFL+uOEVAm0VoAvKRQmnniqT+wkXRILx3Q97bAQPm7UbbekuYQmss
Ei57OA7f49zmYCYJeGALtJPM05TEEl5Q4c1fvVQpOx+YRsZ2ObL3sZnsgRc4Rd6b
EcEEgA3BwSL3vMl1VHqsIBjYlLSUQ+9WsaltSym6sggJrGeMPUxGpbjE/gkV4ltz
wesFdFr/neJNa0RaL0+Ie+gLfNQp1QUHqAF9L7ez89i+fk4q5kv0/0fBBdGY+Uam
k9XEQVZyLWNX0GVLerF3VtRNrmQ/Pg/RWAs9y4x/WCKDD/ZIFFdziEPOL4YWZxbz
PJhU4gGqjY1NywiF2QOLQ6oRN47mT+lb0fYQmrecdRFeDtVdke/gVVy/BtL7zjrd
uIinpcnqUSj0N6Z1NcsRDECI1+AsrmWkQzvplsOdnzUMAAmh0S8KYW4dTixMElaS
1ZKDFAIXjCYhyRi7WocfFSwu3wHGaAQ3UVv1GE1JA6qPDIH4f5wjHK8cBBoJM/Lj
322mA+j+1DwPYbCp46ia1DtMYUyqMn1bLtB6UwAhJr2qEm8pUrdE8+O7FAGIJonm
eIL4aCNXi4gaq1RyiXoAFkayXxL5vpFNljCXGyUG5uzrwl1QFfw/0J86GPOWXjj5
1rdPGzl+q+8vdv4NtWKXjdsLYi3s9LHADnALBi0J6PTKrPI24CLYNrScxEGZXKYf
uyC8FyVFoQuAhToBXZPyxxdQQLw8J7mH3ftMyaya4ka6KhDNMQYuBCHL5GhPAONC
abulB0xuLEBh50rLwVPcwXO2ipFtdaM4EdFKedCKGwk3MuvR4EOY/Mcyx4nPL/cs
yfYwubwJDR7UcXOHD3EORQ2GweeG/0m2ryKNigyb9/Z/9EB3gb3y7AfhaGyiL1Bi
E9e9GQ2sAFUZYWORknN0bYpB2pti0Q3nidBmmN4UzBpPUTpHtbzcNRBc1sylMn4P
pRQebOVQEt9ZJrgq0JGQZPhXSQpXN7DXZwcJk/h7E7eg06p4JgedMGswM5IyZR1J
F9RXcQAEZ/SJirDkg7MRVaShmm/K+AtJOxwN/QFZypsBhc9/PY/LXx0XR2kt+Ev0
IYUbfFHsECFCUy388raxn0d85+6Hy2/JX5EMC6/jFvKT3zWXm4TbxMfqVccCOzi5
bOCJtnwfQIOn93aZuPK/npICjdZDbF62j19YFBJ6iOVWbedsmuwVuYOsz6rZrDdb
K+x1y+SK6gBBPDmvNQfWH+Ks5E9NCPjuR6TG17Xn8yuO9gVys1fTMlGMADgYtWT2
eoVWejeR2e4YduEj6vgdLHIl5kdnNS2gxNidlszdqgf4ln9x9l0UFUbX9EvK7v8J
i4L2sLImCBlfVkQ2O5NgF67Dxp/oeXReRpIaREmI5+VkA4zZMncYSU2g7Yd54cNE
81mBnzl0OZrvUIfCoz6D2361vW+GOOasDAm7/6JstTA03KQmFKK/3VuWFh0mKJ+Z
wkhNcxTq4wS/obQdDAtpBfVjsIzQ50H3ZMXI61p09Qw8NcP5jMFXg+75SnLmfjR6
Tq7xq92f3CIQDWKaoeNsqmiWzF+xDLki6x4O6p0fx5AiLjxamKU8ef1feH2en6hN
BcVD+1zW2viHSM9KUy8zwod/zv9ph97TvzPiYnQ+NJ+myhQwyjFC+5ahQYUyuiom
UZSuI+QGlAb+kLLOXIKDMJ+UtGkocPFAA73GIplch+0DRv7nbhZueQNLL+zVvYrV
gLuaXue8MZQitW4vfpzfx5mEIlNsXQrnMnJx7fkfSl/nFm03aE+CFKKfXy6/o9IW
rYGl5qPE1uVRetQoIXly/uCzF2zm5ONT0ZFl0kBDOXC4yMGQOA6gKlPMsHrQx8NE
ZIaKEzrtpFeoR1x+SnUQad5NsjLUATn49WZJVugaAXLooCJ1/RfdHjuPHsLQA6/b
YzudF1gSLH55RhmfqLNiQfO15P4uiUr4HcFNh3uhGyWezJrL6Eue1jBVz1AXWgtO
V59EXpHQE9T10uYjmwuZaZHc7K+eVH/cvBJlqdj8cKAuZ6Ut1zdzArCO92iccJGq
XDBT7u1/23oTN4Kdz2OJTyJXx5ZDkxil8DOB8/lFDx0bTRfhw+n8SM9dMEbYigN1
rZKq2mGFT0mJPZueR5qp7TMXjHdNSAGvDjcwU7wdd/IwvFX0l140y9VJHgTV7qUo
+eTI34WCYVFJYyGzL2jsfBp9xlsoCaoM1q+u/QVzbBJvGNeoccQR1EoYmZbh1U8b
E6N7SMx8afNqzWpSQcKdRciP0a2uOPiGbYEByDP3eQRhHAgS9E2WF8fBaKKm561+
q0Yuq2kTlzSiuJ/tyNcgM+7F+sMwQjn6w5YuJanOcEZVGQyUDdQHYQOseUvWcUB5
h4v2ueYi1/itnBDQwpQ2h28rEdiX6KX6x8/7GLthvSFuytx4VIM8YP2xJTNxVpZU
XEYphghuYzC5s46zWW8jbbEcCAMNxeALsDhb3kTl0kwZRgIKjYuHSwU6Y6A6ge2Y
yCIGp5B7WiqQ97R58ngiLgUC6aKX6oNwMU/r0RvXg2CGKqI6xSuFewoXgtftVSeB
bosE6T9J7zuYhZxqqJgdEKrIc8EZZqG50z9t5hO346Rv3nC44z6Vti0IK39BQ0lE
3vvhIuFmAHHUl50tbLgzqJ0DJ1NL2suz/e+S0SjDXB3ug1FEtOjRNGyDuvVkrOcr
v4XRJY5ItmJb6uR7q6SGhSxvw+eceFOQSXwDzb0vuMRpKRG7OZJFE6mh1dvtTr8d
jbpCArv43Am59Y10KIGpDeRc89g9hixTJXvF5P5JAnX7KJfwM8Rrp3oWYRv9+jKg
8+MarVGlRzFpZWns/O71Icw4x2bOm+bM4gcbM7Rn+RiElv8Th3KdxDZM9CvGNX4R
dNZyFNPlzLSwF8Ef1yUnw1KVEp5U7GpYv64oOrMDAoC59hCTem+O4u+ZmlCfQPuZ
MmWjhr8AKYwQ5vk9xXh1LS3jbPlWwBw8ra0yof/OOpu+Itu4mwTv6mAA7WZ7efrK
Ua7kD57UFuEhATaZzYnggj2V4p7VPjHqtz6hybGRL/Vf8d/PQNEjpdeNChiihq/o
cH/a9TsTs5SCzSSrwH7HVkKihA9lgi6khIg/vpyLw4bQzLV88lMdbyynL3Cwja0y
yTu/dwlB2GHbhNt7rJ3bM+NY5LOFE2yUvaEFyLZgJsy2DQofIPqtYy5veQP8XOJC
yCe+NEU46uoaFqiNJzIdLJiky+waii2PH/1y9iIp3SUIHYXR3MIi26OS5ciVGOIn
a5zt7CZClyw3xztBi/RIVrpv0uq/Xngf+/z37wX/34raVn/xVl8qM2kfvrK7M6qn
6o5sp0oJl4H5q6RQk1Z7hAGsM1Vr6dlYQa7Z37yovRxxuGeY99Bf6QsvRieR1nRJ
tqP1MgYJN96Dsq94mtF6gRNCqPaMbbEa/P47kZcVR2+De6GgoqSxXK/WibGuvnd3
5SBNpma3+BW1IRhBdTE2y0xXiXvKrc20vE11+5WWQ9QvWDcll+a7n63pLBlqjZxE
fyNOgfBIX+8tRZsJo/DAkepZEHFZkiu6xAuluR2E6OUDBvJZALHO1HISeTJ46geq
a0QPcdruzxX4cQ91P3bZfZHkWLirN82q4ssKB6DSGbdZST/t/jwhzAiqsBfQLLK6
zMOVBWv+/yZ5qG3GWy0jxsBcUmFU92K161hhb6pBZblByBAKdiHMN37xRNFlV7Lb
p/jcsmZRqqwNQlssAjNBrtBLI8zVAPmTne4RSE8pke2gNKIP7kyLFvJipM2Pak5P
FEtlPE13AffxidOVSGBKIdaMPwglWT9Cf94XzF+5xUQjLPr+XoheQD0Y3TXQIgWs
GP02khb9NqmNNTBW+VmaG04yDimYkt16ZXCpbf2Z4XxjQlxMXC4BcnsQeV8F17mg
4VsaTrAmsgOLKPSLKP2r4e7atAL+PaS1tj2E4v+rvc7Z6beVYbPIHxy3aAKxHszc
lqLO10XYL/EIc6pICbD+A+xKFk+IZtLpkVqCJRFzg4Z2laCIQzOgTTPVcvZUdhqP
FxNXfAfWy5IZpR4JhIKlwrwKK5SfCKsrjggl2TlQ8bSzZqYTWknka9iGA7p/kueC
Aa4/h/pZX5cY07odSBTFW1RESy+rgs7teW1W8+u5ogBS2MrnVNHmmITscwY67/oe
CDPAfUimOQC58ANDbDt7aoKDzrI1wPjtYgNfAqcCclEAEYFxKVgkaxuLnr/xLgNs
IVfa05aMwjcRhcWRHSMZKqHn/DkjAfn1EOHuvu+pqiOYI5u9tRAFCcqhFux0L8VU
Xc65Y7qmwRu7ArTMxxJJ0HdO9NqW0S2Ck/TMWx9sOIM62y6hsg6tcq6uogzk2Jyp
0rZHs2omwf6Wkju80T0ouTQWesdfRGEOLpAp+UKOWpFpPAf8vx1n7fHgWnPL/QTI
HvfTohJIaZRr4iL5YmnFv0Gh+EZG9kkmwWHc5afWi9nxRRVQaly6MMe9Tl9c39cT
T7nJ6A5EY4+Ozkwq7k65wLeVi9g9roupWk1/ndyPfCgHNFO6QTH1KGlHYGfGFoML
/CVhleJ0Dwcal695G7+bSl+1bbKkG3kugS9N1iu3Nj8Pyrr4LDijdIuWITXSY/VJ
0ENve/H9Ce6RqrmLcxsEcmPY4QFcbLHkB3QO59HdZkevYSCvtlM3J891MzJhj8Yz
28dO0cjNUOEJYOdeZ/gjw2s4+ZHdmNirfMEiySKhB55q/tQt8E1tNtF1oom3jzO5
DK68AhftA+TGVwnFV9sjvv57QUNo08U2MhbJ4hMX4A2X9I+EJd+eGPqeleFrSjke
LfrZpnI1CHl9OFh9q3lzd0gLJxsVyHpGrdFWC1UB0WBPPGiqEWHhvCpCTPk0Wd57
O20J3iM94DE70gVHv14+CBF9eVTTcIUj2MaA21UiBNSvuAWJ7xKXHcutm5dsB13i
CORlYIRJ/6ENSDRI94Z098BmmjuXh1GUN+8EmREPmOz/q15KzKt319ZiXP8aspn6
41jmW5rvfsK+Cs5GGSGw3QGXKD6g3T7Kud4GAe3uMnicuwOS1gCU0YbDU0pb9Kf3
zN29PR0kesvrBQoqa4FMPQP6gdRj8voopC19usc/VB8K+uuxuJYsBrw9CjDhQbkQ
/6ukdbE+2XB0+0+4uVGIFlHk2DUXEsWYGBlcB8sbQDHrNzde2bsbHyfJ3ZgP6Wgx
Ama2oQg+HqQeNVSV21OY/jGOO6nhWrpsoxlltUzEIRyAA0m4gR0/R4cFUbkdi4gA
wkujIQ494/+VUeSb35KH51a3tJRBwLXDDLPx7tRbFLcuqxspaMGb0QJ3nswQqvP9
MDB3oeN4GtWfZaBYM5Wk2AkhW0f8v1XQs2UVfbvVn/zyYEefaDSG9Vx+40W7fLy5
q9wQMx8gLfC17K8szw9rJDlQ7IzGlYSGL0HShGK16vm5gKAF7eiuRK1clKOj8SgF
eUzoQrIzoQpubz3r3gguz7rc2//FIbq5qOa3oDuV5FbNS43qNkiqKDQfBGiGAoGX
qDTW/R4yyUo+s4bUxEjR2Dw3/peTQfm7XKYBQrf/X/EbhMh/CL/lnhyHhNMqtvYQ
y1CR2k4C6Byn3LAg2uuRNe3KEv3KFlF6K/DJr0o7xbf9Zy+0lk3k5EloVyYfuBYe
Iwbqt/Gq6tTujy/JkXvRWPLoAJ82G+Gj2rgW5ZfUlapy9HAtBrnbpV4ULH6Y3R/r
zh+SF8/CqCSZQcNDz8G2VHIrQzpMAFy5OTcyZn46pHRtn97FBGZrnmtmQhndUmf/
6m0M+V3QA5v/qnrin93OqUFgBLhNm/qLHaOmnzigb1j8KT+nwzmDa9zKQC8iw/lO
ufMadwwtbQ3JNfDu8aLlsry7aCn8nBdubk6C/mbpiU5/7voqNAspAT2yuhpNBZl0
PcqDcoA32j48xVAYgLtrkpbk5xH5m7BsTQdYUK2pL8LIQ8MGycVQJ1fw+XUg6USd
sXvgHveJXN3ElGCoTwElXgNy/eM7UWFGUL9mO1R/+Xf24wCmrJGO9TQ5XFIpQhTY
Rj82iEbctTuiRJCLincgvfyjWcvCzbC1GPDlz870fnIa9eVtAr3/QNCTdBAdCU+c
fyPOgersI0S4SC/6pBi8C2KicsicIGoM7Ire51dDnIMPCQF3PzldrrUelZPk4lC8
rS9SNoCQ8G8KkEQBJdLFJ3ku5r5oc3My2zmreoEZu2tbgTsJWBlCiumfXdpXzNkO
xT73jaVBkY3YiY0ZjLAETXBBKa0FWjq3qloDGoTMcjOX89745k/rvrKeJ0/E5hk2
FYuMRfHF1smFQgrpUy5PUmr0W677TqRSI7p0NS5kIxOjDsj5mhC/CBG+m/LyqDBh
cbJhwuzOw6UsXFAQS/juIcLTlp3/dy0t8X5l6KbbofjF41SYUqlgDQOyX65yfJ2F
lojHqg15b7bZDPKy954dypFzdWqG9Ih66OoJ8jBjUSKo+dGLm41k2+OdszJGzwW/
1TPriyGcEMJV9L9PkDfVtxYxUHAYI9mW/uXMHJq9FYPDlJoI/YPFKf18Ty0eMU5p
YDduLLYoAA83ulxXL9CSohFyF4owc+BcnFo3TK5Fxn3XUHPAD9REjXlTH8QjZkIY
HIBYR48Xz+Z7D53KGSkn3khh0uNjGe6tgT1Q9JkPqruQ4funznSIYkI3F6Q/f8lu
RZsmVxggq/iFfMnnGnBcquXfsO/o/DVNYwgQ8ePVa1Hlo/JLqqJIOfEd48QjwR43
dMO1XUJVPqXaBURquiXY2uDTQR8gdejZgQu3KZ/1Gmfb35fpKdk//Ar3k9ICHvc6
9gCmiCzhs0czOwqKuRsb7gHCa4cKTDsWiEHzPv0fTQpxAJmqrQaormJsRRLAl+qO
FYYUWADjYbljJcZS5/CAjTlExNE2/e+NNONmfIUFLbz9bhYoLToNj3iHa+ZvzkPF
s/m9uIIjUHR7HZ0yeoz2uCQfMH9CXXQugGiG+PwCtMWfIt/vztZuu3W0YiTrPB7x
VfHwg0gMePWhmjnEJIrnHHFjiLIWUQkq7ReGobcDsFxAZ3+8gJHAnnRZ245itQgr
ZU23mgIw3y2qAwl2GnM+Zdarh7KVgL7//2e8bgBU29FSBXknxBgiq6NdW3X38ZH6
oIIQY03VSdeofZxM6ohZGyRKO5gdVq+yCzTjqtcTanBhmWAJnXM2NtUO80e6t8lq
jpJ1Z7oG3mAV5LEtzHSQuGAOGfATs+dhNCV8lpuEJxV6Jsvg0w8TmZpDcVbhyUiX
CSEgu/Hlp9z52mxzD/VzWqo+efWTNQPj7V22Cqj+4UZbXoI17lZfTxIryQKujJtG
rvMkaPPcmw44SCq3DOkpcK5tUeqfZS9To3ykAY2DLiBo/DdX5mED83PU18VOYJRP
tMxVBrxx3eMA52tSCLpcnHoET332ky7iT5a5JvoBQv9iiBUsACo+JxNi+5hKLz0w
MxHWTvmqAPSz9K8mqEQzjiNHdSXCm80cW5/GKJyBwkqdGevZlM92adYLpCaotg1v
l6Xgn4Qw1jUMVTX2x0f5iATySCOoooAhvU69RrYx26y+kF/q/hWqULYcYpo9UWtU
PL7QUbqYpAoVHpVP5dB5pAjFl+duMYyXW0UF5hij4vKDikQ/suW7N5DyytBB9SB0
pmlVFuKYGtAhkFzSvL0F4tj1AkwowKFYHNiKeWkQCb/mIpPDWVo/rKWImFrNlCJR
JSCkuRLnbcfDqDYphjk4VmvAVQh0L5gQKS/Z9dMqDYK2qx6ZN6kJwtrZ8LdE6TwD
1SPRSlfljemVNyMFm+cF3ucvZmuuEbHmnRlXBaFANPUsHKTMkuYNnBwpLsVRdDa9
yP+Yx4+/w1nfotMXCdPlgqb8Pt/U8WhOaotwrmRQzcqB6jm9FTTULlQIeqoyInPZ
kghThv9FC8m1CeJin8EsQK+nwEcNfYY4zrsbxOBP0/wZyzoz/XpRG78gCoRIk77u
HWwJUshrL0mnbCfHR8kix3ynoNVQDYcQxzZld0WQP20S7ZjtTLylvOTnQNhVvGOE
ziJmudz7nkUHzMcX/UdosAsOIHujJoyc2VKUFIJMFXi06qwKWqzHQnODQbEewb4q
NFbaa8St2BKdlaRmNuqLeZZLpsI6w6zM/n578RZGAVbWWbhlV9NRBGCBppMN0GI8
R24ECk1cZ930xMR9A1B2NokDtsAXUZiwQ/BjCLs0PHSJPfvddhYtEY5VWEmRO4sl
OFjoZIz3TfGuHBm6U3fmxf8SKlHQe/srOZENmhXFQpK+htdOm4UzZ+EgHVrcXzSs
iGct5phPDpg7WHrSE5dY1O5gq6YdW/vcva2TNCo44hh4ikr7lLaT+qq2ErfjQKYy
Db54/oq80BKBH2NvSlh8C/ZqWPjDJAFgcCwbjqeFUceOQNNKXhdMjQBI5M4Bnf7i
tE7NMXR78OFi+DYhTGO5ClsqRx30HTcMV36jWeiNAlMxNVI5HIxwYCjpdLxd4Ex4
B80aHDfUtU58JKMMQhzgv5Vxw0aD1zRPjKZe6ujuTqIw1nLkePBwdccCDeE6e+Yz
6o/1snpSVT6lju7HsjrgImGd9z0d9VqLyqBwApjkNKbguapAPCh80Nu8S/IttRHH
q0EizvhLj8e+vEDvlACKC4so12+gcUE2LeOI4oNgIF5e9K0IhJU2TbDkrwVMlCBA
3PD7v7yQ8XDUMsfzUfnMVsRaHxRlFQt5BIHA4uYua90eETpWSfKIpEEIzsG+fcqr
BTD+/9+FlClqhO6CIEXfcNMrvHrdZgfB0uhnRq5DXugXaLK0lg9lUXBFMiQXPHAP
JVtSskLqNM+AIdg4RIXJFa9T8mK00b4EJ641znpp+L690NgtExrFwqSxlDQyATwx
GYyX76pyyz990liIXhFq3m7hO8ypASrvbmEJ8B5b5c5Pb71RvnTU7sLde+EfSS7J
rYI6k0W01jZDMC4Hd+SztwlJ1jPX6Hw3Mxt672Y8MKLBFpZHohJqH4HIraFTXPbF
pErUyuG6DebwPK8nqXFJCE71OQ/eVxiZPrVbHnu97i/9CyqJI0MV+WjhdDE4/95Q
EDR32ugYQQW4/Yd1/nZWRfU0Q/FX/ggUh1rvHCTGUzUyqlb/LrschERJFf0BePgU
394YNBlfhV64i9sH/0ptXZ+dbwMBulBPBStG9lZxdspywm9mBcEAccQ4YPmq4WHp
4YSYxfTXcfM+YG0aoZBJu+oO/wLkXdjiOmOY6rXqIyRkpE9jQq+a+a7JnGVeyCMj
sRUCcmRIboNC2GayKYNvEZ0nB5v9u3VZAR/uJOUrb8CUflnnq+2rbgsVUzAYz9kq
AEY/QLoxGFiSrKuciTlC3GfyX6sS9FDGp5CXA76owXRbC5zt0Qx4YdpVb9MtMs3H
5B/Mp/rsOnuDp6TAzcB8FdDeWnnq5ZTKOP4+F4UFLQsnWXMrDKkSs5b4RUNOoucv
oXG3jv8vWHl2DoJ50i7xzZ4UxfxOJu5JHkBj9JuesqW8dbFl5iCP3s330DY9gcii
uEy2ToQTer2/GOYGn7Wpb8O351++p1ZfCnLxuejyvUOgpIW7xCHj2sBk/OumglC/
sGojDcbz8fjKnDO/p/fENtUw4WDNETPj6rYNHWa0xxBG9xmlNrDgMm80/DdFU4K4
A0DN3Osyuf3FEWIjdkHOkyZG0pifT2lIauQdg3RNXUdkf6Xw1DKb32k5mDyDxcRw
6pE6dBoy6RUVb1GBmzECDcOVgZ/WYI0zks/m9Pvz6ijEuHR7O2UnY/r9jhOMuSFX
FZXwn6wilqHfiX9YkPwPrRgIgzVtmBHBcF7FyNVGYaQS3ePEvrA/VUIUUFt/9lnO
c2wjlbTabaFpUsta2Xku+HuVG4dVoTBcwtRYYYuHuYpBejay890+QMv1EytAIQEC
7zf+m/yll77yH9+79QvXKw/I5zXL67PcO9rnwow+09NBoz8R1cjqpltERmZFE2r9
DI30Y/UxyxdmjUG3SA4jLskVLCQnv2z0FWmI20Fy1SKAJT0YE5K9zZCAMI58x4x0
rvnF4qNAIn9HROSrkGVLDQh6iL0PDlHiFeDYKKUD1s1aaKziePEPk7AoOVtfoLjV
OJTxPQh227Hl+H/kUfEthD3camvpEc9fwH+pUqT2ygtOg92Z9Ke3JFhPSmsBxcfH
n4Hw501i779SrJJAyJFPVembvI/Ay3H3y/49qkLkGby52RApd4a7jzX6wWb0nLNE
T2sYC5KmiDmEWOPddtj8xC7el1spHLb+NNVFqnQrP68scRGYRAm0IopgShyEQFkD
5y8g/opVZGFoRfj6nW0UoG2mWUVXrI7rb9noXSPMDC6VpNzOZ32Q6dz555vba707
ExxU2/A4cfhQaPZiut1yW69iNoo8qG9lph4Ke+7GFGiV41CXt+lRsV5qZm0yS4X4
wH83IEkMdYPMnU5zindJLjyPaBFaugszOrEEWmrKG/3CTLXNjxROX7KPgrmMALjI
mDG93udLisO4tQr21zzZNy3b3TbE21CgObZlwOaYdZPXfUb5Pe+8MnUFd19Z7ryQ
Chmuuuledej++vk4XLifiM9cb5gIJGbUlcQPqsGh92tl/SWj7AyLv0LxS5sVIoW7
ZScT+SEecULTGfaaDE2sbVFIS04YYr8Ygx0TOZCOMl02H2NQU5WphztcXaodYFas
QShocUfyZbGNdXdeMBV7J4Q/z3q8Wm3xmSNwl1fGHGU5bHh4mlTZe2oum600zl9T
fnMyPsJpK2s4w7hQpvYw8ejrh98HDLLB+4m2YgLfBU966jjHmxGnx21qjpsBsOjr
Zxer+aBf/Tol/VXMpD4sM9QSXdFcGItYZaQgjReITPi5j8xhIC9HkPAc0+rERkDU
Z66IZKdMnO853+DZbkFoN6ltBIwUNAYCLugntYcs85OB425N8Fts/mRHH/uDZFtf
QqCJe44ttuktksiBVXEvb6WoVoAoe/TMjqXtQvO0ZmC/5RDN0hjIAmUjU4oGyuLl
stPFwpC/xED/32fB+blNQi9QFgSyhB/hkhAOKiHcOxhipTfyBx5QAiLVggvdguFS
blkad8ldUV/hLfj+SnQNvT7GE0q1nOPUk+2wBUyFDF34OUFS6t3VPRuv59AC7o7u
u4mES5VF0Ht8YdP/X7EC3Sv1zJFiOMLPweNTBQGqLOfqovcpuotVpqtTpDNn3dgp
3uPccEUna1bujubSkvspbYKxZ4IwflzZjWFhgMMDTo9geTVbfArQLEame5uOUzsA
zfQdNpR35cxncHmZofUwh7Wb5DI2gkimMjB17/NRQdZfyDSGasYzAqeDz+WhQUtq
ry5fXtKnKJjEOOqlRAjcVb1m3l0pkUdAcxQiYUtXgitk0Dn9Eyl2Dz0Y7lNl+H3l
ykW2xENertW0PRYDmub/PZH9zdnhXexEL4w3itN1hPgFgiRxChzXq6hT+dEY2OvC
fpyNFBmi0sgZzeoLu4gHGc2EJZYKFW1cumQKpN2uLtV2pnLXdWdEllbQMmTejXle
LZEztlmSVFVIJDhTLOZgbIwNSGezsev8nq4h0kKtMTcHo+ZqLTUlPLKHCbvxc3ts
kZo/l0VlXHul9cW7gDiseLI3/yAjYwwxbQPpCUKYo63bCIhEBvsMAB6wEfmAXVZh
C0Fez6Nc7XKU8sSlthfLPxrv3atYPBfC+amUQ9gj67lgyz1jKWi7fZFYXXc+xVHI
xPT1x3Y3QMDe6LBtB9/NA588X1BdPDUeH8l6vb5yoPksT91mXPkkA05gl/AjtaW0
JVWxnjOvzCkItXLqR1rR4bamjvIu/arm+4RMtzC/assCVnXV5YD+KL8zyzSS0cqx
TgndTEVof+9fc8k+xbxpdG0F8UbDoZLMT85GCY4c/7gzn8ZFosPO9JGS/SqWFxP5
/3/wcMwIqcy5FOA/SlNKd+0BypVxKYFUswk9onC1kH8D7mQCDa+6LUNYvSOMFUyv
A+6LKlDwf3wPzV1qS4567qv3WRwPJD0r6c1tJfCRPukyPaF33Z1pIZ5X3W859o9O
1g6Xu9L+7tKhhgi8516yXG0pPrlHBoDLDLK79sBcKOCqYhHJcOcciF/UuAaYtla5
43GELG6TQr8QHfFdZtrs0iB4r2MZHxg839SdMDKO4SuxDqP7lmgBA4wag8SKFPVq
8Cl3N0LlvgTTziAVqaCazDsc0FfbnfQoOzajD+eOXtkX8NQNn8vaD9x8BPc+5nx2
3Wj5nPUjpqR8QUXASOQV843yr2Hn5UbTtz7Ml0N+eqhxB09Mt3cwam5CzmNUqvd6
3lx7jpLPfo/bbhB3D7B/mzxpHIqb6z8890dOS8p2wPBCLg+oRU8unWK0bIcBk2dk
5rjWBnC92sVYozXbYieI7k2jdQn0BlPoTb36lUxd5UAteFZj3ApEel3OXMuWpYFo
fPPZoB0JWwSI6JLTutCIJY/3Ffyucqb6jzMt7y0jQCIi4NKahhVtQb0i7PYN8Xf/
UISWjpWk29l3WyDOlaVO3Lg9/m+AKTZrHTExaMpCq/bbQGvKeGjKyjBzci7I6vGj
ZCLj1I9DUcXVJBoXFq8VXvUXxhMmMr6k0nTCZITmRYhnCiFAfXVprba2iJe6nj98
n3cOItE1TW1+lJDhLMSws/7rinRBdMcUmECHPdwAzPBhjmYUxncvXV5WBeKtBC7y
6eO2xNyG29WnFXZ1GVKgKZKBNxlurWpgV7L571hXDH53yYbTJjG5hoXaYvp4EUFo
XcyzzzGdIMf0fo0RHLaOl60urttqdYlVM2lN8g1CvwZkWQt3Dw32JR0z2Bylrows
U8zRhdXs4Swsm60mw5ppR1cDorCnCKYczvDE0IomgglHy9PHGhUByfiy+ojjP8vd
5fJ/w09rW2lCe8t8Kyw5Ipv5SL4qRIYCc9vZ+jqSv+tS1g1F+kbfoEtAbFvzJhw+
5p8tbRHXKcfU0Pn7sZvmihu3G0SYYfO2LUDSSr5nqOLKGZlvsKx4SKtLrHUqKOdr
yN7ZZ9GFxfOJ3aILUHD4pyPCiDkipQWuMWbmrKehL3ppO2wSOjmqTE7dZlN2WmIQ
lU0P5AWIEuK9HKD6QLqIZBXz4cgBd7Ur+13XhJX2urRBF+zyMpXl8iwktSDPzIWP
NFlgarSwk2nQ6zP+J++zv+0EHbLmApomqg8XkXwGGlxiFXyck+5Dy1et1ZVQeGxB
OQz2Np2sBpjIzHbOyWX5QNpIoEFV5/TZKfHNT5eCSieh2Y4uTnSCJeeUdl9x4Pzq
CYXEB3ZEj3jwxcNYbv7h0XVPTa3U4n6BtYll3KMF1JDfpFGx4nP0OFTG036zkaWl
NS3qbNGFslrJCvv2qGYz3OxXR29jEZ+7s9cGZl2r47fbNc4cmC4SkX6DWmDmfVDo
QyOh/D1Cl7PStvSDkn7Ex1OWP4XIyF+kcnz/ii3s01TWpJPfML6z8lo+Q0PBiJ1Z
N3b1J8BCRIrh4kRpfcPBQDzo3yeWUCc2YrSgBWS7tYHJXiELI8/er8oYmkNvciyZ
CzJlrCeRCRc/AAMHqzE5Us8Do9iHUBh6cULpjZoZnouvSNVO7tWsi4odek5YvAjE
EO+eRBSDicz92y2cuh7zWGiU3jNZqLUJp6ZdKeJiAy3O5lKS+TCiK5i7EUtL9dq2
ne69yoisKyzZZA3kYD0mBeI1Cj8tZWN4hHnySl4xS/sZUeYVECCymNgD3whHNUV0
eMKR85b1zt750odfLMFgaAPnAGuqdWwg9+gW9GTOhQAGgfLK5h/WczSgSRgMbII+
7T82fA4mrpmOqlxOLY7I0bXztEkBKr2llg4tEz+EoayE9CPYJkxW3mrkGL7KoV9J
r9Y3uQB8+3vaw8h/UJVpHwTceBJZIJFbxCX7A4yRHRzbDnVBhfkK3eM5s7i9qiDp
IQT2wx3+JAhmCVJBAymSMyvvfeWkwrBidJYwKjocIhei6gjELLBrF4VfwJnlsrbf
lQk66uNHM8yePJgLn3HZhMQUmNSFPxsryzEroRcMO4k++oHAFqR5AYxl2tYDMDyB
zC0a62hEuXnn83sQhXUEf1OGGqvpfbRUK19w68YNG2ob/l0EDcB4hRBz63ovlcdV
ge/gIR3FMXlAmFXBmvc7WafekRMUT6r3rwkQKEhjs4gY0osMhdJltyvJfR5VGhJk
JEZrzgqz701o70VCkbxgI7xOyBI1ax8bUSBX+2pVcq2MoNQ+A80pTYi6xhxbPA2K
NuOrQcpoCCFIhejAzmsl28XVF9IZynifOe9DVbZrc5s02nKq+dl+23H8LTX+nBX1
ig1Txk9vwD7Qb0k/OIHdgv/XTKwxge5n/51g+Fs88DEl7NXD/D/TlsRG9m6hUiUC
KCKGXudHEDoGHHviJvDZxaGCo2JgUjaVaBsFRe6MMz1jkj8MyXebso5qjlVZQwt/
2xiZRPvnEESVJhVgKkSRvU2mWpDVqZygd8xyaAV7drj46jtpoNvxabA69eQ2Iwjw
YzF02AJBHG5plmyF7PwuSfFTpkm7nv8N1DqorK3rKcQO/B6MUdra1ZN7bhWF0C3Z
EoOJn3FKQtopNnxT0aDNr55jSWDHop0Lys73c9Aplq48QplgjddD6qSq/hxTxzBy
04m9DzBaPDg6TKA3hCnQW0kBHPsjwrGviQG9ejebz4KucI5xAa0pwp1hRsq8QBZK
MrClwKhH2jbxkwwnO1IRpHeM2N6GkxCfsZpg6dnjXzaXJeUeqIwstn2KJ2XiIIVV
bpn1gPkoEUA1sK6r+r1AwY13hy47nl9gWYlfMSOyBeGBJAEdb60LgWswacSCT907
0LLw6UmnYRYtih2SuBqXS8EWgaD5Yvq2rS8+1LnI/c/UEXaOFbFDp1T8AiNuLLcQ
XUoNYEEfOCuKtfnRGXzZ9/dqXkLcfXSVUYzx9r76kEchkUClAvhpc0YY6rLozVvL
XhC34tJrrSFBOaTJXvRLbcIlYSi7NWPISpiIvOQcg4M6YJHHzl/+FL85iCOZu8tq
Qi6CyauvIEKQ4wSei+sKjMFv6AYqh1poPFXfCvkiPV72cF5alJFIj2GjQl/i3FXq
0Bi5BqOtHzNQ1oD6jb2nJF3FLlTfNDghDqV7mD7S1vDkKtBPjNvsK3VLhUs5bTq7
5PyiNDe7fzRk9HD+r96mtV4SGjsr1opjXwDs94RpMOJ79wlVNmDo5UpgJXG2PA6n
08tYVRnkLxxTrJfphwkhUxYaZjwx8lbKyIztdsiIemzNnGy5HLpfz0wWTPN2EFFD
US1okIqpQdh+PbaH9gVw5c4+Z6PUJ/0LeNuJgBLTxS6dxOa3k7OPoPS2rIca+Ycv
JHD7M2SAAN+2KuyR5721vx62SUOBo3NqN6x4rVRHnmARdLIUv+7g7Lfx4N7+vd0x
8f5DrtSZsp7YKTRKZMQ5fLAYdOW4Pi9A2OFOmBf2RJ+owcxV4FQkhxzAziHrDh2m
QpVzPOOFHt2jnDcOVvytzU81P1JQ6K7c4gXjoQDeOBJtackn90hdBYG0Jibaed22
rW8n6bDLuq11tc2bCu8rH7GJDMmYSpIagMumqQ/dOj8JHF2Kp9JFV4CZEv26Wb/U
1ENjtnO2RI2WYRkdMZWwgFYK3TCM2K0R9LPcQ2/SKqIPGYfMmfcRYjqM5UMIruin
HPhc0nUYfhMM4A8YdThu63kLUBQbyvIjhurDtzncggAnRJMpszA6Mziv9Q8YAt4Q
/dVTbduRTUOJg5Da5eBTrY+glD+Ra7k2aD9EWZFZ3yYdp4YHST6uQSiG4yU7AOqr
OIwT3ExjjnIvuMJ3vu4aIfiGGdxyKhxdremwr6JC3wTOLHzX2lOVA7qCx0sY9xPM
MDfCEVgkCU1y2CtsbeUgzsAtqyrmZ67wducClJEDm/PTuoTYBWVM17nHBZ4Sqnft
7Al7ZaQOFFuJoL6TmnBO07Aif0+aUzqxuchXfyIIiyh4OwZLOvyCvO5ZibeO9jsI
rtyMMADELWg0mNlUyh1RClVinVyPPNc/bKd/zBJ1k/rUbylzNCxxccyMMwBciL/J
qwFNZRIW3RTG/iXEHJ6x6XdcZ8N35myVQqzD6eG3rZrwL9mU31Slm3O8szCZXDK9
B3e4eObiGXP9NyGfkVc1cj5jR6KZ52G3+KzyQlorel9LXjGIOc+kPkDAI9gj0zIN
lttOca8lrXBgCa03fhVHzjyHQC3fgayn3FAreT0OLvTXioPMwIZKp15hLUUx4pBf
n4FuWf0JfNoFHKP0ZsdC3To83MEU7hG2JvHvurSfXzjXSX6yTEBb0RAQcZ743pQP
WiUpP2A73NwwsTVk9J5CjkHDY7qvdbWKfGQEr54I5M/CvPUvvtuSR3JEZyzxgSq+
dgZJ4vPFzDI3i/I06P+VXd8EtGBMSni+X4AILqkZKuK6GRuSuZOu3tUxpMq4MYgM
3nrhyBmBeWUcdO+MyKVGP9QH3qKJeCFMSw9uj+PPD7P01wbrtGJoQ+eHNG1Wad5y
CAuwDZY//wLp7gkHgscZepkrX8jS8rgJpp2fLwhnw/sxRZfxT4PunclbCrznpnGK
XEWWhquRNJB4iSpVpAkS1r7TEHIhduYstZ1+ympp7OOJ0MVP4dcYuLF+7/n2FnPg
OwpZ0y6dC/YevhQDROyxMW8IWQvzgaA+3LxkLeu0vLEYttFVC/02Y80tEPu4D5/B
lAoQ0U41gdLss94nCM1+F2w42UFvF9tCOQPPGS8xKgnY55I8TCY/R0h+uQbbIFK/
TM1vi2xdg7q2a9V/DTtBvM2JBjG8jKQVJrxOnDS2AiajiEGxrFDp8E6TRL0g9mv8
vyppf8JJSwlEFs0/PYbxbRyiKNZn0kUDOugIabXtFxWpmmO0Qe+BEBqGBmuDw4hX
5P0bVIFV6i52MnQ/iovSFxVj1pmKX8+qCuphLAHfKyz9Up40/11t8+ckochJxFw9
Kec/Tmg7ubwJwEqFRA2Hvh0t7yL8dB7EpTDF5x8zQOoK8Ja5eN4uLE04+PnzECVI
2kZW/u0q3zzl9+TF2dcl4rjsih4z+3o+EpcGMMaPzGwEwpL7I2R2ULx8E3irBzp/
ZGs99+2dgsTzo6zqNtzVN4jn9WkiYUeajvoHLMM1iEAgH4arAL8FrakT6fa83Kkx
79eaQZe+yo1jiUMFnwL+NHmIZooo/Dz/tT7X08NuJ5oem36VRM9E9oy8G1fT6gEy
Ap3mWxKqON1TvMX99FTSHlEqa+Dv8CrBMaXobILNJTSTtYj56c3ms884X/dH/6Rq
Au4GwhJUZbUjhHQVtLljTVtJzpI2Lnd6CsLKB8Kla3AVtlT+KI0mcrZGFErzn2hU
oMCBUwcaSjVlA9pLoJtvAnWt8D47QSxJfNzqfcoUbC8ssjmicC3gEHaPvdypyuHt
3crYNv99WpQ77gXViMqO7gi0B2uWqFFhIEX8R4GDhRiPXX6SGwak8OsVxBN+T+VL
QXyApYao3NaNXeSrqzpT85HpDIi6rpgUc1vnLE0nWtg1mmKKr9jXx6ccW63DQZJE
3UJo01XunR52FaBiskRcr0SvmrcKQ7mQMvsga2+PqfVi0hsM0tKZ+QVHYZc8ZAs4
bNbeUPUeEaJxLkiAQeinTuuAAOPpmpW5bmddpEwPOPw6764t35wRbB0nY4zLVQDJ
3cauKTiaWZXQRfMQJ4MT/AtLekVST/PS736YLGmVXd4JFDMU5YzmN9kAJLIZa93p
odWS2HEt9bu3i2Xvx7B3NQudfBxhL1/0/v7vHIN8jE+QD/SgP/JvmsoS/aSNORby
ADu/NcfeCnkIf33FMifbJyEJwB1kJ4SXJRzsWIkbUFj+/A7TurWqi6Uo/lWzIrGH
FmaQvN5L6KJjcE1GqheyYcNRHXE8NC3TztnVKqmU3Zlu2yB1yhMxewRHWFvwT22N
U4eB5fnQt7u4yoXwp2JHBy/CdlBt50kqqxK3cq3sTzUrufbPlGdzPu0hAxq2A/K6
QicT15gyPsCALLCCsIx3Y+0duEcoaD4UPq8MOKxOtJrsvnkJx3kRu/isEwi7UgtS
HVVSvs4oafGTMuj7/FFQOon4LtJj6Fhvr0/QwkoLOF3iAFQp6w++8Io5bsy1gl9h
GkRByAX6nVrm59AwdqRPGHwjPQ1AwXMdnS7U/6bLNk0oEz7RH7O8IZlCFE5WPqPK
sWjHEXNix3t+oDKoqVG9OtsGrTsuim3CA8fsUZVwp2uW3+ySN/2QMo4/sUVna4e9
yeacbKSFTiBFS8hvBb3VyqnNEzBdb1wW8Q4VBlkAo4AJR40aFjOgCeM+jFf+VOU3
gIMqOJx69xvUdT1J325bXvNuK2+3jwDrN1FbJcDQzGjdj2eK/mDg8eIQSozfjCVS
nSKx7OKQBvr5sk8YGcOR64cqwUCUU5JGoUmvlCW7J6wQ8oxLoM0G7krbRBFAja51
JJA2ddBODLlv1pS+cDzUJO/3oY64XyYqVaMdw0iygpGwAZRJjghGrFQTzXAZs9e4
btp4wMY2F0/fSYAtdsA4XC0IlKKMBnDXSLLCWFTvN7XzpCvxxh4rtacbAF7x0VDV
BARauv4XsV4HRhQEi3ofFUh5+7cdLSVi1NgTUSO3lfe/JEyjlE4qSioeVHRZxO22
29/Uv2bgwqPPMMXkMHD5wszVcYuxuERCI7NF0YH9BgIHbgLK8W03Q/PYgxXe2+nV
ls771VVs+drYJO/2U6dxqhMLkukiBGPGOJPWIvxCFP1ynDUVQemjzvcd0LLNhzN7
zqURfsIqthfcwIkVqlCK+9jTJxpC20+XyoVxYMG++fFQ6dzDoGmNaYa71mwgibvQ
ZE15bBevsrj6Kkmf/WQ9CpAJc6Or/w848tpe/o/5DHBrBCFK3Mha0u7NbwFhFS8I
Y6LLO96i/drq9P99VbLf52TWwUIQkXlGnBIrvA7H1yOWsPT/4j/tKwDbn2OqHhZx
REH5leelqnym2JkawhY12+ghubfRXR1eocd7bMY0uiTXqLurKNKzwELR/52S6Aop
45qEYWcp5sB1GYSCaMyQ43+nnX//xrMXqVQonCwVYU40w1Hs3yQE8SXCi+HGZaW1
Y+SIFUb4trbSoro6oZaC9svKvI1yU3qoAArPS426fmcjfdFpexEUtAyi3nR2g2uA
04GKIgJFHLLbCH1SrTkRXwmu1kVNan3STFVBKByUfAdE4EzGrR0tp2UumYPTL8kG
lM4FbUxwii0JVAcVD6WU+Uo2aPhMqAPFQo+xb4OpqKL1CF7l/4tZjv9Ti1MzUwoL
XoxEf5rQNFO6060E6+tg68/CNCi/MvkZ/gW8wsy/71G5M7ahMEyRQQBbNQA8t/Je
B9ls4ItrpcCj8eSFPDe/MzkHXKkUredKpQaFrwqLHrVNY4xBBieO4V6yLVggxVF/
zbBCdupZef8Ri0YqqJ0u00s77GTQ4Y1+GLMuhro7Hed4ISTtsg9YSdHxSPjQ/iw7
i79NZbf1o2BwH+Yj8MbrQE4ijlOHV/TdoaMRWYy+Cnrdgb3Q6/UubR3tNBTYkIsM
KEvUI2F3Kzxjx+aXWIxnRL/v3XoSD7OVMQepMopeAZxJ8zNPURckrEAvMYHoP6Gd
Ty9RmlN2zDdiKwozzxngLJ252I5liSoLA5TmEq24QaAe77P+IKxu9/FYgCJ3BBAf
EljbWO/6OiQsYbHX6qt35fJMj2XReZhftJSEHUh6/S3n6Ovf9kn0osL0/GD2reTw
fj0X9uAPSP1FBvJyzJKNHEVPkZp0eV0mEkKsYk+Y42S5dGI5lYmxQ5BbzZ6cJHJc
rT7yGsdxxkc5XnaFVeS7Uhdb4X6cmnt+JpW5T6jbd53yUJ55VwJAZvkHDZ3w3nZ1
DUXAJK3MhyIN8lMo7vYsSQjnXY+j0aiOFqJR4MiaXThVVLhYAr87kBMK1jgho3Yy
sLjmRYe00QgNqD/sVhU+UC/+UluttGVCisA+Pb6MOyYPsZHY5aOenLg1/1t2G8wS
u1/H+Xja0HWQKu93sUchkWa6vzhHscOjU4idWxKr7oL+ojvGjogH2vGLqehljYBG
0R3XndX9GWGecLq+1pAhORM3ezPOJiqssdVF5hb7B7KUCHQW/ABdUGY9oNVneNR9
iwM94BtTKtGMEV3wepwgGJhORjsN5Hy0A2VcpQSQ4TfHMo7zWr3QiLspb2Xt9Y1J
fTigbPwsfcZ0D7BnlhcRv2AO5slItF0JjZ+fIvdevTN6SvRu70Ri1e+EFwSQqxlW
nUvKIv1vPAojsxq2+aZWf245gGNgkuN1amIdWTtK5LBCja6JBehHBChRIeFnNNSX
3rvLR5cm9H2+96iLUCFfIu9r9t4Xnsr3A61rduRE5z+H8bYEJG8FEVsqi+G0uGwr
HdUrTzJ5Kf4nk6pBVB5cTHK47XOnQigm6UUFg8gfko9UKeQUk+sok6n6OMyI8w7h
hhbBqF5/mzmew//3C8rfsN842ydeODW488ARUIoQtWrSGp7FHgsTtxK1K+rZgbZW
lyUKO4w3VGUGILUcbrtNelJ7FtC0Kvup553DNDFlWfhW7s0m01uS4cA10FCz2rkv
nInpud6cqDms2mPkzdbkiXIgWgKXlW0gdfg8fdeoISAGb+AQ+IaKIbapUQrKlmts
l277jN2MXdVuir/lP5bKe4mJB5ZW80skejt1QkbIlheUwOM1yzhfFEVjrnld1Zm1
8qSFZj+YHPIfwNRnXJY4Tc0XRy8gX4cFjdzSQUf0cn959PCkgNjEUUMdWkJzTJJC
vREkWwg6JQ9rHvHDS0q03gP3aEoNWSu/ZUN3tc5FfSEkhH5X/mjRFffFduDCmKVW
OnNACR42ML9VaKluYxb/IhMgJk2sFOOa92MRcR2EpQmU58N/Udqcis/4s5kVa4Ip
GAsF/eMus6FoJgcsl3xbCRv8e2x9NDkCh2RIVaHah0GXDSSbuMI2as608AXw5PPe
9tO2NcVzXgp35kfOIj/ysioB7z243b2mnXlNLrYOgBOzJv3dawBGyJyIsuLyCa+k
1gvDoG939MrDM1LWyFguvK6TWanIojB7qsyoSqZQ7BNxykAo7GnT4Cy3YfaMhinQ
bgxx5n42q8hQkMWCxPWgkgbM26ugRyS09y8oEvi5trncdA1uEDNBX3AEY36iUkU2
pA5woE5+IkiDRYmHz4Y9KiDdOJRKcmr2pHssUerwUJlC02ySvAtGu5smpUM4kCP0
uoBHIes0BGnk33tbyhfDMiDyNFinCb4vqBp9SVt2e9EXvb29pSnalXQGOyepf2Qp
CMX/xVIG7YgdbExkIMbgT6qFBv8+i5YvD/PTHjB51EGXlsFHFzkoSHU6W0ifhCSC
UvA8ACf5zMEmjVmnkzEI8M6Zi45ap7soB1L918bthTlptCdUQcMMd4HcBmg29PcY
8OC1u4wsM0j754MFClMZmrKnBUamlWzosD1XUWed6cve21E2q/AyWROdBw8ED7RU
+3Z6Rwu+V1D2kyrMlUl+oXJQcniNa5xlD5cYlXAtgYc5D9RWbDDQo7qwjXVKaq62
dSeyrY+jK+LDYlrfvbypzkb+PuFwyz9jhsHTH5E4zJuAqtjxMo2Rdtjqh9oEBgo/
3oI1hdslRKywvlhhV+6HrmpoEG13W3kR1w4cWDlWaql+Qb2KJqFaOzMXlNKqhqRQ
+zNIOEp7Y9vakaglY+h8kryn8qK9nWgms9jkLSzESUS1XoHRCWh06axzY18EfH1n
iqJ6zF8O0CTIsoSAL5hv3vxaS/mXoZaluQnupUFzgeuRm+ey+n0S1iQIJZ3TEQEN
bUlLb4CSJndJUTe5ek0cY+YQ2mImZgqXV1MJO5JTxIOytY9bLqKiwvKnJxf4rfPx
tpHIILsl09OtVVHplm+JYaCxLwIqGAw2tnkIVkGR4dFjyo0fJ+iwSTDrTIJbSd/Q
3KJhk8/797sfUTTjH1D1WrU5ER2mX5mofa7K3in14a4KDPIXAkQlNDJH324gDN2t
wSmGAQczeriwpvc33ZYpxfqsHuyM5I2s2OMB/YH7ILJ6XkAsnmraDlobPjBjt1QY
e7JpqX2tBPIjrFoUmfXC6WSAevE5qlDK43enzyb9gOOXXdNG22+4ihF0G5Hm0+iE
kGZ2+ayH8NV4q9LBbZXWdL1KX96cIsKxO/fM1bj8k09SZdtCl5JX5XZ3E46aTTE+
lbM0+U3uQnLW29Xc0qa57O3YOmeugdKCpjBfy38QzU3U2ADQoLeyrMSpwdEvyC9F
FjQ2GCvzpLta0sxRkcOsKp1KZ6pe3aYPME4dLN6Ptqi8CJfIbjBil0BB/zBFPjfs
K8O5sKaO1vL/5UxzFdsN4/raxJgzPYU1EZwka/GUO+MLZZj7atnJcxCy0hbCcu/y
r084cIaSOym4FunNfLVHov95VR6j+rCw48PVsTqGWU6LDyxkEComcS6XZ+qEPLMG
K9XsZrZh3GMwINbmSzEwoccFMLCXMXFLSCtLYPtWT815ewucxPv4i+f98MLjaT2M
IwAXGh8gaSHp7liR6E6OxjV62UfKqe5rnppgQ4cwNg0LJmxD70BkJErXXhmmDxW2
8MNC3Sq4X25kv0OY98D5x6DeGF6PA+DJgrDOaRenNDVa67IC3U/3LFVORlciDw+9
cjLIRBy4Rlvwh/o5hpAhb11FEDAu8MWA6LEt3vWGBlNWG52QXDH+y6jck6ZgSat1
4/CWpvkGKlgjD9EekfVQ33enLX+gdG3kwbYjQcsivauQbXe3CzkHWLTmRER9XsI/
hGKtmwj22ops2gDCN+tf9XhxEFdzOv6Kxfa6l4VbeOW5wCFPk2HD+AQGomecoyL2
A8e2XCCbIOKKslkjkx6EcmsjFP8uA3YTzSRV+6UomDtevTlr5jU2zwNOZwwlKAjS
yrY4opRGgaiVHsh/qhCWbjKnQ9ykQF7BfbvaVn8YzMKijbhL6iJlRzXbU/nsXznX
nEyLiCTCPcArKn1DoPhftXjb25rTY/AWEMKH8/1Tly1ej0ahSiIXhYfVOKVA2vIj
4DAxXsBoX4GB6kxrqnUfuYv1U2s9ZtUx0qb1MOp3g8NKBhUWqO57aBTqEiTbkOPX
rZJD2I6eXkIKHLLIJsbeMI0tnDbme3LagnNiyEiNljbH8Jz7TddOkXMGaISA6vv1
qqFIvQuIqV48DSQxYsqoAyc+/TCIqfqxg7FBbr6itXNbhP4R7BJeWocgfS3+xeUm
LgNsUeXT7JNaS0k+onDe8R46Im1ZS4oLwsBoVERjqx2UnWebfvyLcPY8P9BczA/O
7GdkGyUt6k2/dvmXWUOdRAE/sM4rfIVOwjL83uNH4HATlq9+JJhLTOSVlRJBUspU
Af5R7s8iMvsPMlEqWB3rDSXotsYCEWV10kS5ygW+25FXT/QcTca11qgi5y+aoV/g
aTB1FVGAt/T01ctXEMzUrKhpP/VALItfH/hNm93YwP70gTZ1Zy35MnoE6XYsYtOv
wtRw2p67uFbk8reM1UMW5qzXWY89JzdGIkLfWBCgTTN1Wu9U9+gXaJIr1sKFiUOW
cz8NHcxucFPXENf4LBQE0Ztcy2GgaLzZCHc+XwLjQSklLtqhwUGwVTVLNpYGLNQD
zK/DgAcDgxBHINeTO5pFUtuI092oQwzY4rs5E+7oZjnhroD4JwZUsYk1W5/oDM2Z
M6AObULYz+PGlnoFbGmirR6wGYQ1T95bPR0deI/VEgvHBkaaYIMPekOjVUsrali7
ZTDB2ONHbX3XgvrMsSHDRlc9pmk6ksxEy6dDKug8mpBOVmuqA9fzQu/WwyVtwSOW
WhZv6H5FtnBWD0tz77zsagWdflwZY7BVdPcTrEkje9P+WH6ql7SE93fS92KBXfh+
G1dT22Gg4jviIkxAFP9O8Qb/A54w+0PBE5MuS0/d8Tw3L4IYMbvRoi0o3HqYqNSu
FLL3wXcQR27r7pdtUuLM4YcnOyojsFny0ChD7+P4HDWkut85tIgb49BlaUqKuRzL
0ZjjedApBlxeiGeGuRG8zpk/qqYVi1Q7SzkO/0p8PsOjKlt1QhHFgA21wWjNCxPK
gRwl7YwXSuMfzyZ6l+I8zzUNtyJJckIEfuiVnX/prvPi6NBsq6j3m0dLmzvgfH0o
eHSpR5AdJioqVjKhWQcpZH2h2Y/D5STm9pht9c9FvWkg7IniHzBDEcGYagNjJ/3K
m+2g/bPAc3RnbA4IxXfV6g2g/P5ITZhMHGSLhcjXKrs1l/pJpe4lZQJrolnQ1nCR
AFHIPH3si5Ttv5DLqU+p6xrFummDOHkoseyKDO4P0agN581PBarNjq9XANahur75
6erzkyB98tECePz+dG4eNM3bJ6aVpCNkuUdnR0qBIlaCSF/QE+qAchE4CeJVIR9N
xQdaagXSEr2Y4eGQhe/uRrj1b5S/kHxObBeCY+OsnwOFrFcJKwPskCe6SdNdJ70c
cFM5NdzKJlR8sNJH3tPaKoFcFZ5RKwIHDZgJMIqlNhyPhq0paaTEyyaConSdQ53E
+vsLOCE8JTlx3iGIM3jygGmXjr3phh2qs1j5+nJYMpLyHeLJeCensAQQmulfwdHm
KX3UDJrD91yLgdycEBnfVwWrxph7f2+EAuSKI1hJ9/POIcnwsMm/jyTBMCeFpaF6
HQLkVBEwgOqpRLa0IvyAKb8FcUQnnh7cjv3Lpctiz7CY4Uwdm+B8Qx3RlWMdOZcb
9a+COt1wwBM0yP0xhzVOT8Gyi0E0navbrj/DXk0wG6K8kRtulGkttIzs28AEwXBi
xES6bg4Tb/zkREQTm1lp5jfsUpQ3ioeRybQspbBLqc8/fP12mjGdLBgif7xPa+fJ
8vrgu/uKnkGrRU9SRACHrbbRQK9vP871ak5T5Y323ei/tIZ9KC5tZdhCWRs0KENJ
GPdnAcmD1N6dtAqXQEcJnilP53pWs6ghU+lGcLKJPK60MiNkTQPG8dp0W5PklTHu
Wjp1NAzbFrNv8cic6TWEfm2DsMbEM/71gzk+HASzgW2SU78Q3pEH8+L8vkVD+rVP
qKc/YQbDheyH0wie6DP2hd4IGMdcZ67VhvmKui7IF0Ij+6Ul/4F33Oo0oDcOrcE4
5B13Xt+sYrF2xhIbrnYmwOHTtDOheUKmJj22mvL6iMGvO5XO9ZBpLPO8WTLI8zK7
54F1KRv0LdSHdjPtIFrmqQT7y+89GOmRj6YOfMvA9yjmJr+lngt9Zi4hU4L6rW/p
IRLBr8idHFNpbfUuc+hq2/SHH6cjb7MgR7NbX8ZAxXdJJLLJb/oNQ0afhEk7+Q7f
PJu2/MttVuKf9oBHsbOitsxvChOJrY5rhmK7u+Y/idMQrw3UX2V8Opd1AXr/NGNn
Z8hlmTKTmgmrat2/gM1G+lidgb2BbtwCEDtCMkCuYrYj+OpGZE40/Ct0OOrmEhm1
4PGxRHt+jV6ss2V7DdSDVfB6SeIQ8C6AUVSMegPvP996G6xjuTjBYTUgOqvkBxfP
ehsNJ9lqvfDzlQZrKKffMCHj+77F6NPiVXTEul+JkC4jUZewHkQnOoaX8kpdzdVz
RUYKrlDgUeu4ekymeN53QUtQUrDi78Yr+Ye4+puqm9Un3+6jYFpy+1RIM7bPW6uq
26qEvE2/z6ylief9aPhUQglynx1oQCIlL0mfk/SrtAhvQoj0voQGWYxwu5Lzp6oy
igsI+m0y8NiTwcsqtdr7H/q6CSO2heilnyVjsAgrrdnxfoTqnwYxVMt52PQt9oUP
i9l0DydLbTbTto8AQ9yQTj3ttWTMgRY/2HFkwICYSJSE3OAbCIHeRTgRD3DznnAl
L5djDmTHAMCuFwz4KK1UCedSMgozHfzwctYg09e1FIpjCondaB4LPY0CBFTLD1Uu
/GHUS1yi+8WC0+TV2eivLbWToW7QRZqGV4QKw/Ur5Ziz8l6Yrzz6tZYb1fUw18cy
lJIuOvakpWCqwncpz8GJ7LEkwFsU2eIf7tRWltp1Y19/u/JeK8F7D1vUWDHcdmJU
FJu4RuEN1D0+puMrmri5g1DTdYboXi6HorwDcveZpXc5a7J9o8OwOeRzT1oVfwJ2
zUPCFS3vpZHTKcLZKTScKBBGZSq4ivmSQqPBatm7394qh0nY43zVZZwz7oITGtsu
nB6tfeUFP+W5lrFhpgIpeeigt4jCuzJd9+0Ayh09caLmRk4vCw+tP3ZqA5Y9fH6f
wADFNLtNXRPQUZYThQKyK4lZH/5mPpBr5b4lnBMoLEmnjZG9p4kx/1PWypmMM0F2
Tc3Y6NXbbunFC1ScpFGTuU52Z825v878dEfHNcUSNFgdvK+Vqc3ucOqOowEWLxmd
ZPSDI2pexIXjA9OXNaJQkG/N5IcLbxR2XwuKeDiGw80cJ/wU12dw4VlTec+L8Qrc
syeJsiUX/hb89XQUbxai16RXD977XG0sj0vMO4mOn8jMr4cCSU1YwzEzPVxidcq6
RXPoRxf8POJ9KgVO92TP5RzTwudTQigg4ipPZuoOesJh0/fpm++gam6eUQ6+L5uR
8lE8sX2zWO6nhuQWrh2ZVc863Rij4s5y42+b5lH+kVTKpv1iRqGN59Ikr2z8D7gD
O0plCNthygZVYmdvfvHtug9EDenQFT1yEVANukz+5YVONZQj/QjmVKg5g6aUkt91
auDnqm0GSjqUmGsNlStdD/plFZrZWd0WJBo313cWnvcxbqGFG48qidmAuVtqMAmo
9cUpcbCK124q92Zpmq4Sgb40nCb9IZYiCdIAtFa6znPeQp0lGM4B7ntTDsEz+UD2
Yqg0IWSfH8qUFwgry+0i2ANSNjgJ4nqNygO8HDRwV4xdAyq/b6Hyt1xnHmYcfcvr
43nWDHnD3PbrooAEGBeYLC/vecHcRbiqKP0ARpD1DdHlwsBcZ+APUSV4paE4xDGa
WBl1ihYGv196docwdcsL10jo/vGjGLxlNi6h+5WVMEf960nF/P/KJNDKdfIIKGno
k/C6arNvJl1O5q8Ub0NtvTjrhZ0UETuZOU7HEUeEP9tITzfV8Mrw3lf+JqGvs6mc
pZ12akLZ/etHSCMpg7wYXGaoDoXPA0B2ZLf60RHoZNBR4YAPRKzVScJQynK83ujS
dFgBRoFDIkFZGT/qyhPEAnAgDMTaRm8gFcdxNhNkPPD1z/xKO3yDLZQz09yx/p9U
NEeU+9wyD52FCGJk9AyRYL/9nAprGqHJg2BM7QWvUUnEot3Ch9Em4Q2ckTQ0DHxB
QcoVX4wx78yPkq2oyOZWtdl6aHhtOxoTrWFjicfNJtOrXEtymdmoOv4oWocYXFJa
FmbkAsR5UR2UGfpl10Su1HVRT2DKfX/R8mJRUJA47StwhTUKPWhavl3m/GrtDtXl
0bDGFOrLPUmwhapAsQavqJXiebpFFBYZip5/I18IlGprFd58AN6DCkr8B+K1+JdB
Udwky/O7ruCaWVASc6vDlboURPJQxR1SFJfV1z/McBCeQmrtlSMPMfFD+Jkhe/oa
yJaS9pQJeI8odbHHa4+Ohbpstkle45Wd8IkxbY5/5+ZYDfvC1TYQmNtzlUU87ncC
A+pWqV1J4HLGg7tMwfhbVKc5p8UFeQ08QI1uDgPxxDEv51mqnFUkSbBkrvrCwaF0
02kunntZ6Uy+J3Uc6K4jT6LH4uZatSR4o4Bvz1wWe4dPD+g/CkI887AwIdEn5qDI
MW0dGy3t22nK1Huh0ZTE/G4dA/ZWiUlTrnz22JxQhaWTQF1ZudJ/tNMlKo/1/msU
f10A+d1X7zkDH/+kfhd9yWTJiShj6WB18dzXrP0A/VIwgZfkgSzzHYDR/ejycLGE
BiHOU58EHlfIfBAGLu+wjPByW7U2ZXzKzfr7QyClsOskSIx7gXY3kHU8SeCc9bH/
DW/AA80N+jPnh67yAHccBT2jw+wAxJdaZoGXzgz3O4/kSqYBaouSwwPrawHT68xl
yo+NQTrPkf6E3mp4G/MNfqt4H8SFVggiBSEFfOmWbzID0Y0cgCmXDklhfD3mW3DS
0A7js5IqNnWKiGlS8NJh9hmtfBsXqpoGJIUCWaCND7nfQaT7bdGkg+IHRnqw2h3G
ivGIBXyNCNFxch3l/Lf/aritf3+ITjLX+mTPUBywVltecd1o+POrh1jD/Lq3u49Q
LLyftvrPx7n/kyHvWqhMZVWO2gJr/DwLAwUSMyc0PCd5DS5GAMRS+6wy2bZh+spf
vwDhz7bgGvyPJVJyyvL/W+sDrMkZfZUqqkEpTOcZuKYdvCLQiGWyrtUSldetvxFE
2DxUvCLDuvQaxpbZdfvoWxXfRdw3G7ZFzfEpIrsSn6aYYbtkQUHVlz3TYmXmzAV2
Wvr2mJiny1bUDDMqoOCsGkd+s4bu2Bk9/CqahJwtQ/AjT/qtTGAcTAcvGSYeTjLs
a1rB/s+4oVBRmeE0PSvZcZGb7NwOKpVwqwkpjaXydRUTypLuRtCirRqjzAZUzgiL
9zTUN5OmWhxmfyywMq6DMUYIZqN8pqwXf7E9iNBQXf6RIY8dkZ9OFWadQWIVZFJj
yKkUckDsIUkNIl8jT8GRjseArVaGqlSvmfygQOtps4T6s8JuOFiY+m2vZskZBzee
xw8GieOCiQYjPcJuwr5ItcdIbzh9jSJAqi9jPvrFMFUDxqMlfAz+74d8mhkVj94g
ky6EBmCyCvK1JXvaXRNNerFd6rU+1Bp42P/S4AAGY0fgkCJbEy59zwxuO5b/9HhC
5DqqnuXEBLSjqIObqa64rvZ5JzOets6FR0RykSL/lqWn2XSM/f8+MkjqgeTN1ase
5rmKkhMqNNahlxaD4jHDukac/GDIXx+4dWMnnVq8GZXlZNID4tUnfI3X4hGr45Us
p4haM6d72T2YIsBr+E4hkW7kU7K/YgcegCLnnQqZS5nEmLsvylyM2VqOFHtQkiyH
6zhgA7NDfNurEmffFUB+HsmktLwPxBlwesJc7K4MsFI0OzyeAju9v3lg7oUTZxfQ
GqYs9r9LSh+Z3SvEnXE/T1DTdRNfWX7lvcxhz4hfi2JfjWNXIf6r52wmftLaMtLZ
qUgYSYIfq93q27R7MdPyRa7R25N5+dIODHF6oC0GY+h8B8NO9+8NGTxgOiDmAmG+
a4mwmV5Y/KJnvuDvRkJQy2FtRsVeEo38poSAFKq9vYDWjq1MJFEiUAZ7Hz+ZilxA
jLT8hK+sUiGFzgPmL31ubVPXJkHIWqwiTeCcxlx+9NMlVoxuUwVj6NdbXgCT5446
T9+IwVFX0Vnmi+KPvqW8E69l2iXOV2HUGi98N6AlfifA2jryRMVX5cPd0BqxLomX
vj/u4f1wolRvxKOojyo5PQkgYxnAREvmcJGlLojeKKo7Ijycp5+DEl+ZlWkOWr/7
yQaTvnLNu2xS4P9nRvwrY4SMA/SbyK2FpKsqtIchBNWLUY8AE3D87o3A9AsQ44CV
UYkHSNuJWJ7rYNJyaYlF53mYYeqnAtQ94BNPOq5alh5/vC0qEsHArqML19M2A8KP
S6188Gk3FfisJj5rG5hHQT9pAO2EBSTpZEYfEntyYA2HIRLpqxpn/weKWqY+UTAR
xvNyBRZ/Y/pVa7Jo4in5WcYUODQFU6ypPD5j0gsLBJmTztcYWGiIDwvtUinLThNH
tZC0ImdaNJiB8Ix2OVQ54SK74O/BIrby1oATnABM2ZTfOcEtYvV4jBIhKIyRE7G7
Ks7aoJyHiRtmJxgF0/TU6mXGKAXiq1EueockOc7GNGhUhuHjMeKu36IlByKi7oGG
glcHVBlCg3iGq2U9Q07gt4nHeTaSTCnI3gWTL5CMLREs0XsPakt7OqjFHM7+N06+
bXmYA7vVJHkPuCQdB7VqMg1wHLpUM/aaSLxgSIo02yRiqt6M83+NKvZy5SdgPzb4
X1oJZLxtTQBZ1clAZGdFXMlaR8Y/zW/h+yjasCdgxVYhR9Xkp1AKxmNrRv45Q9+0
IcgT2iGRXii98taa9VLiuhI5jBYjEceUv5IFZ9wz+I0t1cCnf25ULcLZwKj0fMwk
k6XCXrR0mx/VHsgt4Fcj0DVXPPoy3+iMkQxaGtLezS2c4LjvbScSaEMJqrsVc3eH
jAG2PsUkDCzTb0LWElpB9YfwbHPg7gKUIh1R1/dT07faAgrtTZRGgCkW/Z+vszhA
Nlkq1YgFqINkG0z+/YYh3uIrDgSg3JHQ+mOkfRU5ajCVUFrIlB8CROA9L9qFFFJR
woGG4Tyxj9ub7Nd4YWTmq6yob8EHQ+I/cD8SUM2sRZg92ECvzA7b4Vd0C42PyznT
qLGad3XGP4CUtfeMoeo6bG8AKrtnZoVznBaE62QivXh/Nl7Fg8EbICHjbLgosMgN
yf6DP4MUGjFHjsq2C/dtBZrdzo6KQFBhqSE5bLzTuLNHbB8Q+pFAaPJmkw/G/feY
/IgOh4fHhxAeXP+IRhwHbMrYqUpsWqXkq/8oO94Xknq1p32bylsNblP9mN5obsBz
v3EShHKqP4Db41tGCVDlldh2t0xFaPigJazgbYwhcEAZSLhwVwrYsvLz3iXGhUVy
AZP/bm17BArFh/4k/jW7+wacpoZacF3uHLALcLSQE0/+enoVlALSgjPylLORuzLS
ySfsIpOx4CjBYKgmRutg8nvKeZNEU2VLsW/lw9aAp8+GmauyVdh5i7PKUWSiKQOu
L8uqkH74hdMsTbr32zXE6NXEuDxfb8bULqR7lKjXPeZtHRYsvlU5zzesl2zT62aE
4Fem2QSO05J9WauWPL8vozbUGy6TWJ6UBmKNzEF4F1neGsTALkqUIrsUjA0VmYTN
a0tR0rwm40yqf4Zwhz/VhcJTHjU+UQpfDKE6kTXFTaQyHn79tk9EAHUUCVVMp/Pt
Vz3orMN371sNMAh6mmIn2eHWHR9xO1NUUsp87piBgpDoN1eKEnpN1nUQjBxE9JM8
Hhgavxg1Rpk8plA0tIGWZw38hn6RC70egMkcneIu0J679TansfgNvMEIxI2unU5J
pYr/f7fGQZ/BS8qQsQ+qDL+FayAwjLtxOEqYd/ffLl/Nx899E9wX+RRm7E+0HKYX
5e46GycdHhMHnupfGfrBNIncoLlt3wdCtc7zyyZqx0JgcNoyNkIPSSTUsAj4gswV
uzGo+PgWusNFNOA/wIVnVutc8dspwEvSNcev4fTRGi4YmvJWasnNtvkA4Qu89bPp
hBLLn8LPJkiQ5GhuF5riUrZ75b8BvPO7e22j6/nUJAY3B2UIqEu6Zt9O5pYBVUNH
KTYD3Z+NgCiKTieAzVhGADxEWjDmQxVWJO7hG0+/pSSnw6iGBP0r3Lam+R3J4Vv/
2fyj/p1JvoLjuu7BBGGU4m/n8erLzqQH5odjhGh0hbD47gyPn3JecB3LElTM6T9x
X5EYM2MdRaMGZnh3ZU/EXhooeVXDJIU3EqQK17jIjnwSmXeDS9CTJfnMoqTFBH39
7fA4p+FO7VzshbGug4WrfEj18aZ/FONF338XTchKFK4yNEeu/KsFHpNCeo3uAd2q
qmhb+0DlxfhDLPrk5S5j/o/8USVBrm6Mn1XxWd0zPE5YjZTfbCXg1Fe56Pvh9ydj
QTsEaX90hyUcy1IfOzRYriEO1Fzvr84fBhIlz/3BsdKcgJLTV00sBP/QdXkI63Zl
GkLz6MY9Cu0jiZwvsq02DkwtIVCCKqKat5p6oanQHMRrIJa+rC7393AxZYMzfdoz
wfz09+4enLndiY3Kjs67Fu3yxM925r0UlIK20c2FDtbPNqgWV6MaI+bx0ISQYEHy
3qHTadcmFWaNGiU/9uf8wIyfwCohtjhHSflpBF5P2Kq8YRgaPILYQWnkg+EQcX2C
NHqcq+1QHWvxkba4tfbXmYe7RKjXqCsrUN5lgNecM7pZ+Li64B88FYz17ComIWZL
gzo6YbXbUNoM3kE6qTStP+DZCd17oQ/5Zz+g+bSg6IASQKKI8Fglpqd9diaf8lVi
MTMref7GBZXTeO5UsgxiHJpEr0FQPWpWOqNMochIw+CTwMRq8l99PG6Uv4jJqAhP
TInpRvif7k0spUqOCz5j+Pvo1QVGqikAgmYgzVj4EZz0qfIh233hw4V8HM+31xnx
G8hecsiA3Z4nFbOktHRJGd8FGRPI3jcJksd2PvC0XijhUE1M/frIf7MzmJvaZ/d9
jL6IwqBxSCh4z+RPihROTbZ3pmemHa383d1EdKhCBu1J0/utl/brsKK8zaMIWxl2
1wKSjcSdk8Ss9wtfwBcs7adOKVUwpL3CJalHDtVmJv0xe+Zlokz7LrCQIp0rKeLM
eprGcb/aM1XEh+od2dH6DsWBXCVI+rRft9kTkXpXuj0DeDJoMVeiSQCLuqHuL+Pg
C38B+rPe5BW5m/IONeM5Mlvz99VYKI2p5FWg47TSGnO9GyFe+PWwHXAX92AcrXZG
OT0WiGVYJqiNkcIUD88d7/hPky9N6J23q1rdTt7Zsv7gbs8zHqX/rgCfGwbUs9GC
GhyVBQCsQFV554LYPeqdxOQxe2Rk3+vmSeJ5BWFD7YXmTV5A7VpxlD9I1YYYm004
CQSMdmap8RxoZPr+7F1dg87R8b0WOwxFJqYYv9KK5oRSWckDb9SAx0yA/xRdPWH2
TMCpEHUqFWIJ72SZ0VeJ7m8HHSNtcqZYWjst/F9gcqcj+zR+y1yxH6HwnHUQ02dC
yCkz0+wVkwcSOP0Pqj0o+xSDrsBBvSdjOIIHRG+BiZnq5JaWij21JU/KXxYSXWZM
CZ6XIxtVgAxgIwopPB2x2yMyXnZ/0XG47+sdEpgHP3O023U6FU7GLc1UJz8lM/Mk
L0Cc/ByY4cw5m7/hlx/NQ41LAz0aPeoGNs6Qr+mkrnI0uUC9Y0fbvrMQnd1Uhe8P
S67g2c4BKRyuYIFBzHI+uE2xebxcRsbJgDRqr70+KZOE8eymMCGrKkGlwn14VB6A
i2Mz9qAmDc2qBAK8SqdXWVa/K5ASGB+tYly/4c1CbCdD8FgnXAWL+f7vdf4fdccx
RGVxNSDogTkCK/AcY1d+xPMMp8Ezj5M2nF68fzc1SyXbxV8n6gG9vQxDGzMAi4ps
drtI8zuEMszsGWbiiNd8z4+wItxW9zhqeZXrPE5HbVVDyRlohcnZUZba3VUxH8xh
a7cxirt9F9xWB+EPCYIquUxm8n0lWgu5neFUSokcEo3IMsrd7GUqeWNjHsga1Sbg
h7bzmGliZa8W/TDhatoicmFlGDboX0ZHG5RuXwHdTpO2O6/E2uFw5ZfcXpyXF9ky
vGYSAsDEjVlBb4ZDUg+AEB1GHzw7Usq1zmqC30YUqJ37lBH+pIc4waQHxopySYYA
mQZinAIL8uB31ZMie48tI3zxX5pBXKN8o/PHEUL00q90lt70FnQpW46o4+VfqGRO
79nRq8l/q5HLXQTZbkQBAjW++wsHLXc18PL+DWvSe2DPvwjKTX/ankXMTZjUnz2i
kvPW+fitORUGvIQa0ky6FV2pTrzYTMPPsGry+slxSfWyyv2Ri5CviE9XlbfLpM68
G5+UX9zQSeL9cG7ACk1R9ALcthovQvGXY2As1KqFNnGntcwNWSyJgj6uGr3dxqet
VV3z16bF9byJhuQ1GrzLSTNGHGg9gNhyM3ScAAVPzymvsam1ab5iawrFXzdfAisR
9RMlk5NQrIfiPXau2Ko2pWiwKe7+Ys6vkEt7GlWQlpO4y9KWeQgQelX+A6qF5+Js
Y7XU+xmor+0u1X2ebU1Wd67N/OzEN1+q3Y6/nfFSWVylNfqNX6at+nM6+DJuYrNk
oxxKIQJOMFuJKlAZbebx5KyaWUSPt7gDgzAseRDOBdg5Jyf1ehiVBBgDx2BA7R7/
0mbjXk9xTTTlNjWGd3bI5LKjxqMDPxqKCca9lRHK3++Er4YgN8l4kJ3J45nGY3H2
GAMky7zmsmYMOH1YQYppgWQL2JCp7AvgECX/If3ztQq170lFEZi5BRxz1qkeqOyb
DB7MbSsvzkKkNJc3CckyUaXdto/kwa0gEoKSHN7OoEiGoqACfBsi03STbOimHnEu
LzscIWtl4AAj5HaSQvL2GSspxiMHJ45KqtL23/nBBbuDTEneUKHgS6urQk8Thf3A
dhQ02Ar8OMDRzsERuuohlp9DoXup9u2X0QOaD4gg4ACkha33X9mGcWrOhQbiEJel
zUZ1YAK0xKIVpaSm7Y8Ow6Tjd4a+51k1mBaSkOUdnB++J3eAOX6QwaXIG9m4LO+K
dljk50kMFGcsM5qvGnweERY5wlbmEkDbfptQmN95ik2yCZtZeM+ytBYQHotqtSqc
i/x4uS16D4mToTFZZl5XNSBJvpsR313ovXsifLtKZ0DbQOMSvX1fAKgyk1PRxfyW
8kgiitakPRdzHUFlhj5OEB1PbmtjTLLOGDlBkrv2TW7oiJFJfKBmG5a41eTUBKRt
89htCf1wIeLrqaEX7G17OCCWwSRFi2cUPkiai/ytlrz6NUVNzgingY2600XEVYUq
2AyhfNvDF1TIF+O4a8yPVZfNOaOAh0VgExGo23CP+WNAnzInPBTVKc/PGkxGemHI
TWHSP+LzE4DDGUnHSpyVnlPU8PV8FfYyYXegc49+ieYB4xI1b5ni6iqx4kPIHlSD
m674de9pKjEkD6GqPsDMaGbsdtHLlS4Glb5wS06qarRPAbe3kzYrlXP5mycPjldm
sjR5LirrI68CXi1mx9PzwwSaaiuzSTNVLss4RivrjZ0hDoM2Ksh4OkBjZvyLOg0v
fx/c3z2oiTVB/F0CGyE9VJl3RYvG7n5F9IHimAo+nwaVDPGdD9Go6ZRuJV8xAQ5Y
Q7J3EXLoaAFse6OGdfhXI0XGuyPqCCxNZmNHd3CSR3qbA5i89SXrEjWOyBLsUeHR
QFNw77qRxt/PSkPl8pz8jKe2dTVVHuaS4S2TrWXh8cSWGQMqvHuqBCib+yKZixLV
jm0dy6jzjQRW0FByic11eZeq0xll3aAP/IdBbJRCzkQ64QjB0cUc7VrS5FF/aAGt
UZzSYyxgG0OxDBbv76Qk0zlPrG7a3VS1K/o2a4CVdQ76qIL87I0s/3kM0bt/eMpr
N3xVAgdwoRGS4f1/cQkuuMLCX5T4SmK/5OJz0+ko47IsB/MqR4KwaATI4lRn7al5
naRHAJPigaCvh5WGbn/rpgeceCPag2xW/ujz9BPG2VudhmjDr2iFOO9O8Hk4yL0X
t9hr4ljFekfDAfNS7nFjsz7EjGFbd3L7eznf47UY2mttWnxQ1MPmtHKGBjETZKGy
knjMBnwtBQsy9KpyZ7ZSiCNwx9gkNWSmC+G3Oi8IinhF6mzhVzAQyCWeDUkJDS4R
xDUHWMQcYwJPbttugO/wiFBOMANfitXreSrxQT/OfHl2krmlpOeW90PqzHFPqWD6
7I+p08IatOKnAkpl/dSHQTJWP/DiVhwQUddgzT2lDyY6Ejklh/JN3B9nTbTReThR
gZbAYf3h4OnjggUUk05niDZBSo5HJxktvTffuOuQ7cXvxYr6XoMmoxYcCBJrIlXO
ZsDxBNXb82d5gixVDJ9uOgeaxUBPs11lSr7usA2k/3TsoHVFc3KQO5gkF0lKfFLm
yR7Y3LYkRac++as9K+2WLHjs+x2SqGzDrAGi8l2tiLM/tYfEZooVVVVk0OLr0JSA
2fQdvJpCBcry+6B/YqbS6GnXnoNqLinxC+rEfL0XCML6yBqIfTf4ZR3RCPF+Z2H6
SHM2sIiVregB8O/22Hu66Pn4gHx8iH4ZMr756aBYhgL798CmCQIQoDbKxw1uoPAW
5PnLN/yhabtE8O5kLHLsRBj/Sjmksyq+iVV12MVZ2Kt2yn4h914lXdIlzVR89/1Z
7YrXTM78Qyrlf60ECuXghKie85jKcJb7IRIfvg16Joi+VRKimGrpQqhE2STQampX
4h/CwjUgVhb1qSPn5F0kUIyDFG1DaqKow+8x3pjCcdiN8UwReKzS2isbyQHzQHOt
i7wLYAvhnkoYoD4v3lNsuEP3Fbn83EH2gNigBMbeQIysc73guCdlPrFwcg1AOu6g
wHDg2GVWpNDHk2n6lmDZ9GuY20baP/ZkPdOE0r9RxjtCVJCq6aBCtYwEPid8I4He
ZalCOOm5ZKcmviVHLDgfpR+mdY+NiEaznf9b2kvf6AM9jP2wT/zfBLpL/uhPvx94
jbnxeV6AXMKPMEQhKD5sUK5ekTy8IKxWWn73+6b38KHL9AckFNv4lmBF+RxQFfzs
Lz+lmvZ/H2xI7Kj6cS3OJBI6Ve31v0HQHror7Yuk0KyNdrkd0gt1PNOJd5PMLosP
a+NnAlX7w6KbWe+p4XkUQ56Nc0ujX2SnTe6eoKN08qB3l2W/iPKLxzy5RVz9BfDH
ExGnKYikaUl3Jpcfh0Eof92+VjezvXKV90/lCrir8tKdnJvm59UcmBGvhdvXqs7f
LQTmQTPxSX1XO/YjRliVQis5VRubG3BkVEgJTbsJCB8R39eGVaeCbwAO5R4RgQTs
J2MK8mZu+OyHcJfcRvR4HZ0p3OVZ5iOUFV4vVfSwRjoprEhk+V+eCpLMxuuxyGrg
aHKFobPpqL0ymdluPopTls9QRh+S0AfuploYHRBAk2H9b4NBVV7sZ96oU6oY/JfG
yJIJ2fPAnPMsQFXaYYo9PlwpuVsgSzb7y0p+WYDJYCBkQW+L2pC7L4l00qVk/aNb
QdZg0iG6DJeEkhnq99VZw3MXiRrEVS4TpGwZ5+b7kATYHvsHbkIEJ1O8/PVCT5ns
xTrZQ5QyY7VXxGYnmlZ9i1pKjipX74eIXl2/KWyqSO2vO9JtpJ7lqWwzeCa44OQL
WR+JZbXFUXlOkl+L0pG8IJGFUZGbzG8nTk1V6B/GVFtOJB9o6K1+U3o5ATyL/xUI
MO0t6bUuWF/JJWPQcqvbVrUhYtnt62LE4EsJhacCbBEpEpIioxIz5HOeef+vcicg
E0qr1UVPgCfec2oLcd3m/RdzOx7KPC+Qjz+lTj42WgvikyPw4YO2jgGBIn550Lbh
Po9PhH2P+HKbtHtXzlpPUAtUZsMLxY7LTic2g1kh/JEmBgQSovXEkZefKNUGaJrZ
mqzKQczOFop93/Ts/EnhJuisabruYF2YTS3bZ5lgMD+4j2+m6Zi/7BXxh7S+/egr
++/yIQwzVesGcsay95aOIYQttcaNNBX/i+aa2HgJ2ZBrw/Sv9Jy4Tns0Sy5SDqGI
KQ3KKX13qy8NQEX8zUyGMXw6PP9SnzmJKLJWnsM+Hw/1kPG4gldxPrtvGx1TlAvp
lsyt3vKlhy5sk5/VOPKn50vddNdQSh0FTlNfjcbwMBzeIBHV4lTza37VwNqIS2Gb
H6NWYeThnCDgp+ChKBzNQ/cX9o26RxjypHWclyzYIKlo466Anv1keQ0xlP+dQhIJ
/IpgY5DR4rgKc9ws21FXuDaEJYT6qzoCk2hBeU8gMVzXMMJaO22KJYBYENVPJ7yV
9oeofkT6bXrlZ3rG6w2g6dYShdWa/bj45QaoH5A6Qx3joIwaNl4yVJRq41UnSP0q
rOWdtpl/RIxo/YJKo5HG7GOTQr9z0dWkz1ALvqukaNvTCJv63Nk0nUsUO2lqBXgK
JZtjkVuM0XCfG5XLHKUyzYMTFGnLTGsKYoLJHGxKzE0y0T+1flr6Ca3UbhtNQCCf
gIrWlwWLOhr+LL98EdrXYb02FViqpEefdgvQQhrX2kfU7iMpNQ8SMw2wi8ifBm6p
Csn6ui4/+mzKGruuQm3Ls/p0LqmkSe9Q8i6RwXnZ94yPTxX4ZZUEBFLtHaUtl77S
EDhAT0LZzjYO6oSoRHfpFFRrDZEwm+PBtU+enZut9HEogJW8tf9rAV1FLSZr/U1e
Z+MSIC9x4m/yMLt/D7fTAAGycRipzcrN0m3egBKraxfeBJ99AxPKBSOfAOgahQEr
IiUmZgysjeWbOTNYa7LlkA7xWBtnEn6l4p/v1Geu8ZON44s2hkn2tUzKzf63bs9C
9bAPN8Fv2c/46j5ZRlYLCdYyj6cay6O9bJSQ/qSBlKLoqM2yrt8OjqEOrMdG6NAK
wynhduUakxuloCrwG0XhTUhE0nxbh1TVI/By2GswCO43FKqn6mrY+KkKimOs2oa+
SyAKbRJHfJRxrqeI1FMUQut/ADb8DpxGLQ2QT8Fv6SYQNeuvepyswUc+wr38lq12
gzbtTSxIEStn1z63zL1o/hfR8Bngb0KgI+P5ToxuSTtBd77LYVrrxYiAoaFZEHM6
oUK0tcPhw+S/O2NDVq9VLQjXeJqfk4HC/3yuCsuQaDFUnuZlIEvcLAolSc+2jj7b
IddQz+XS6OttdcI5Six0aXIu5qV2a1Chh7u4kvc7OJ3669RQpn19qoaij7F+nO7A
tHVERQsoCbwMMoe0PlFhmW5IaSo328mvypOIomjAJbE3bagWaUy2c6U5JdkUocwm
j4soEksoZNZXHOfs/wM/2kTY6TwauIJZFPbiStxiwde+h2VnVO4vvwPH3nFrXCqD
ksSCL1xfauGbFjpFo4IzbE2KiYA++5LEEL3HSESQ3bI87op7FfEX+uvHBUk7f4nC
SLActN2vrqt/Gn6IObHHfLjgJiT2CFNVVwaFOo8cqwtMlGNCeVfmzPzrs/Jv1Teh
WEqXHaoZTPdi60Ci/OKLhpOFnXb6fl5xcgeWlGUKvDL2R3YdwL6Gvqm1MtVU9dUi
a0dyac8vaC2cHq34caCl3GqY8DjSkGa/x26B9mDliC7gLlnIXh1nyrFF7A46n6ki
EIPD02MiYyi14FfHwgMuR4aNjt3SZv/jonl2Y+ZqTSKTk52D3FOccPr271iH1yD0
6L9diUUbL+jlNpnpNI7gBweyTyQSCIFQbQyUmTdTOxNN/xZr3zl0/hI3AEXWJDL3
VlvhqFjuAtTlRVXTnoRheWCe+7TnrefmXANZieJsRzEjOESl7nZeXQtf6fzdiWjJ
DerTZ9IiQ/ux/gWXAU0VeYxzEZplmRN7xZzHIINhJ4tsW37uBmcPVRf3ZH5ILG3P
ntiYQ0mtrIoa0n3syLypJiIgvbciulAr7r6aAARyGiMdYr6CVKyzlDORGyvV7O2M
43XTCIrV1bOxVVCkrCs909L11eAwcDItwRvpt4pFc6GFn1KjZl4yADJliqZIQgtt
jtEW7nINLkayEysAGmIDpWR0rXWl1PGCj35Pe1eQ93m3ilTA9i0nqR8T63LIJipk
pcuv84usd5v46QPGmC+u2S7rRo+LKD784EMOmkeZMwqgFlldadWk9+Vc4MsVqBBZ
rb5DxOEyXF50dkZe2SGfRlvhj+bXQ+obE/EW2wQZhXRPZH5FoRs82Zjhbke55Ryk
YH3TPQ10TT1TPBvzFW1b3KGNUbrtsowR7NoxDSJR7OjSEaAElCJ1Cq9OAMyyR0Xc
nwP0+ruKqoJ0S4tiDIZSUluGOSCJlZoAOf7qrIbFWGaDtLkPoNqkeWrgCo+vmW0G
Q3mfZp457WccXHhQOUlij3wExLUSUU3Fl6dqmXvDHI+iDbiJKXWox7U+5FUAWRKM
hY0gphCEJdN6eE7PiD78gi0qvz0MANYhKo65bqdsrvtRRQF0pEoeYMGslbYTgqQT
iJMXGFwaXF8erGzRmKY5jqhuYD/5BO18Hfv0OaIe7qGU0Ytg2S4aMGOlgO/Zziur
TNsdaAcPYUMwcyM5VdRsfHohJ4bF7hwjsOsaaJsFQ6SkFPlOVAGyYtb3JrKMh39c
ckvY8S0QNw6+ABrJlCPxteS2+XnDkuaCVsfn9IlfCYb+7bZMnS8E21UEqslNOhSY
CxH9WRk7PSm0C/7CveH2/KAvc603jrff/Mgq26BVEfm7Z2XcZStBwc/qOI4Cro17
VNfGTb0P//sakH+rdyqmT/be406hgq8+lOPEJ0L7Ju//Iy3SbdA7g4Fv66R3ekbz
J/B013QFXMES+RBN0n68YA3eJ2GcjOYIhPfLrROxGjc7sPZ9prR671OAA3Dw2is+
RXr+PHqtUQe+bK/HNcfAQaXNNaeqL0ZDobMhUG0mvVeDenqH74hS5ANPYFlv7svM
2tEFfG1Mf2ulKrOjx9tgqlNgJ5L0bh+xuIsZVStnAUqCSpbI+AAFnGIffwF0p6Wp
H8ziA+NUZFKQljsSH/VMvRKzHX2upym+lRhCQQqyXuWamL+yYTNRH26TJf1kAuHr
Ez3g2KXfC2qHDm/86JTyooD6vsqaU6wlBE64QA2z7/HpO4NE0Ul6JoLdyJY3zlwp
zU0TBZMo5Fid9pHLQ9Z+zfDnUfvrIEd/TwGhOfA6GBVqnq14BwvvVgmgz3x74/tX
g9Yw8VpR35jykOIsJTNIN/fiov8nSyFKkukvYv5qdasZB2fVcarf/T96+wLckyHX
DD5TPIO/TPiTRRZpJA/Yeht756cktsGmFSKyzPC8K+BPFyxnRlBrXCpIe0cFy0jG
o/C7dvjvNJqqgCG0Acn7dV38u5U4zGy/sNikdsbtYTEvQosOMiImxcWY3gTtNa/f
d6zHFzpp/y1YcFyMFrme8uF2K7jMQdl8BmNzGAmpsajHgh9X5j1f5wfHIYPbpLgS
AyB4rDLHzQxSsf6R0yTVA4L10aYhw3GjYpRN4CQWgKVrJP5G7q06sqt7PjPLSRye
rt34vFayFYH/McHTAAwRWIgKGSuSJ3NxTzc5YrHSMHL6EY2RuF/s71OsJfdF1h81
iVRYrip+Bzr2Z6LCxL2pC6gzUrt0DldJC8n8VVtP9iMAG2dk2LRQzhiUd2cQDbxO
bDF7puGVDXAaGlO51QEAANWiCP/OqIYhmFk77zgkPLokyMV5VYcPrpCAb5pp2NEU
afPpprF8sEl4S/+upbogpSXUaLH6XXeYtBJHQGfsU0NidOZB/LbJHucuyDszmE/3
RZVtnORKBS0oJuLWIab6LFZB7cbtNaZjaxJbcnEuxxS6NAcX6uR0C9kbJTy5qe5T
zcG6eeUntS6epQQRY6F/ANyHH1W8ND/5RvlTijiZXQUzpoRxrU67WXNugayxG2Wj
VOWTHjh2srSydlxGZnNw6Aihx3GtlcQE6EbDGcWqikT5iCiQoqZ+e2pCYvA7n+kl
vcOeWy/TMkNoE9jUyTfnIjHqA6M+T08rLmhLgeYw+uqhWj83/Ad06JEqMsmUGURs
NTg03hKD+Dz3SSRVouiXhn/WlffzquLlVMGg3IeG22fJZDS1kouKYtUqNZ8s4uqp
jeEEVPa2k2MgjOGc91tlxv8JGP9MGP0zNtd28+XrWX0X51kK/ox9hYWpgLTvThlM
Eq1mplPotUsv48EpkMi9QfisAbj2Ir5ppERQFFA6Et+BBb7By2TwGjzOEfsckwKt
doIuT9UY7Mz8sMiHVuFUuyiPKvBksZfN7eU6NNlUafxZC2HYq2PEZVNubLFV0ttQ
TV9FVOuKMspsOr7v7bJAnLmZXpifa5HaNc7js+78pnDqyvQs8DBia93dPr9esBwZ
rHTsZf/BrKcrwpNTkqEN6hrhzrpdaMvSZJA+kgtHlCTZ4rkuj2XwSQY+npEPKYwU
zcNOJtTTO+JKZNUwa/o+3VHFFxdaxNeuJNCcj57kCz/wl22xOuSRZnX9Q8cVio6e
OumrK4dT6fvObwMH7dqibBcP+GRthqAVolgRnCb8AAmERsmKpC+NtPKU6st2Kkuy
x9nhaynQJHeyCTXRPAVu7Bb80hZmyJC3Vv+ub0HG59lnZ5TUYLGFbYExCez/g4+l
5UL7ncnon4MnVrdQ0RBqV8CGh4vIVjEvFbeYUYV09Yt8QvQcHwDAC7+f89lBTTgo
GaTu2ZGzh4/STakF7iX8/M2y4aOgjPdWBS/PX/75UB58NQXO0JzoyQzT9YiO++f+
JJnKAgUwxgH6Oce2FndEfelwOz7zxtzL/tZe8Q7oMltINzb0IVqLl2m4mNk64BQt
MC3bT5PJUyrzoG4BWWD8BVdNSXjTLZgtgNxwK0CU35popy4zLKFQxQXTyFuV4jyt
U05WsDQ6qSUxc1zN+YmpW08GsRdos529uu8B9uYUfavxutMUtnX4o087cPUsWkPM
ty/iQo6aid/JDg6UcHv+xIQVCvJPHlsjlSXoFHH/T5apLIw6V1TPVi+OQrUOhZn5
E869HkgvaV/awwNHNdDA2GGpENNhaL+ebhPejD8P7Ee3xIPeDi8hxSbylQxny3Uj
ajCmB1R8d3GwxzZH0R6eH0Cj430koRAezIrItj0UQ5hvnnBBAd4vLicp0c+3hgvz
vObffx4w9sjGZzEcnneG4Np25m9anDGYivS8v8wIHf6C854sMJrX6BoosoOBJ46c
iHu47yJePRDfRs9+IDe9cXrKezThhz9PadUNkJf7bpXuLyyDudE5pOTpmQ/Dw5va
pHEvImS8qy+HpDazDy3dRvLFfmLPUEwN1TBc6nSpTpQ9LAhq6cI9lUJQ0BXfksfR
/MiCbcsTeTQMTTRc84yh9lQRroQeCZLcVyPj4QycvOBfr89ZTLUanHf+IeMn8rUX
MCJoT7KWQ7WBbj3Nii1+fsdPulNjBzxwd72s/EGug47T5q6qEv6F630QLFwLnVTy
Cu9iHaNm9lwM6jKdl0hKyspdX0+fx5jqVrpcP6QYv4cPYXtjN0wKPvlukQI9JObR
S0JJV2XTTAJjuOt0R/S5ri+zLHgmmhgVRvrwHYr6/C+xx4Rt0auYEEag0HCS09ln
KYvx8Zg8PbkHIcIS8trHuRoHQ0qKQxfqzoK0NRM+Db/FJPY7qAFQFM/aZy+8RsG6
5izI2+n7wIcYG6DWbmIeOCU1NYKsXV0ieaBtRQXSsmc7Qdwd+eukcVkGz4yE+Lu5
YHOnRBNFfJMUYVJJOGZbouc0jcUJtYPzGbjjYzomhOD1LEU2c8dnS7SI985qC+Lm
oL4otsOS0yhjgcAVmrvOOZ8bZXIAlL+tBS+zVdLPXM0BZF1E6U1kKJX240XwmBZv
pGiGxzMKQk7Oh1UzyveCmC3OY6YDXKlDmo6EcwqGbT35vtkdJ7VXVDFPhLeecudV
Z4ijC8njL8jiYz+qGSyfn2ATBx3mvvY2gGsQ9B2H4/lU2X8Lbm4YWZpWQ66fmp72
wCqVsp2chQucphmKkhfrGtYo1HKkokzK3oEQph/CX6mOf9fOlHsTv9cmbdR17SAf
BbPvcxTGzGe63EFKEMvTqIH2Ohc+grVShA8xBIJR7FPy6HT1yqL79/JjLIJP9pKX
WUaoHsBx/LLxGUeYzx/C2vU+Omb3+7xg/A3PZsnB0/kGMzE0NTgemNHRztpEtvmS
eKo6pzYZ+fcHxLC7yRZmHB2HZKHfdhSSwJfv1vcn7JuaqLhFo+BGg3KQGog6XdRQ
ac/mADCgYnwnkaciwMX4hm+GKEjfUGCUFi1lczOvkANKWJIIRAEdYamYzxTnGob9
BuAOi/+ALO4i7M7uvNN0Thh6jPnaqwJQRFWmPxQue58ryXvPoNeuMr8vn/9Nvulo
Q+oJRx1SP2uNuUZkcyNoYd+JXFGQ/YkNnqfGuxYkegm1m6iWG+2ZZFQmhPYmuW8g
DG2Q3vmcpRZkeHMAAydR8cZIkT7rV9nRiqrJ4LHkNaoRnDPJyJgDUNUjwj3P/Ovw
Nw0N8n/QwG0QKiU4yc8pe9fRDbHi51eVujqWQC4rGM75hxLrkcnznKPWkcUWNUxV
nxDFPQxClBgoNqy9zCC5D2A+Ev2GkIDXjSzUzpeQCIW95lDyVX9+WdXqc2xfH9QJ
VtWXFVAAZ6FAwzN+pepxNgmhIUK8lS3kh7PbfcFCHxEd5usTGfjImDZoxT8l6UaH
rTcU2btHY8KwhA74oOnViI8lPxFrgy41Js4O3fSFzw6tIgbV5gmBKMrxlcch71qC
XvfZLNfDKleaFrn7zAMGGbxMTi7k3iWEz3E8CUzbqN3JOTbfHfWg7S3YFMdAcLxl
3Tq1bS/ppRSYclOt39fKPVdTML+4ie4gxRakX8iIqYmxjlSux7MS7OQ3eOzB4u3m
kI0teBNByDgmHqQrf4ItUYtnJRZmdH/yg3LHPK5Jep4pjjAom542y0ma+2kh8blM
0eJNJLTM/k4fx4dSrUR5SIS59f4Ge2xZQwzF+FKGjbmrE3AooDgQEWrP8ZCGZGHR
x9lW4+l2mmYnYV0zlglanlYI2KrWtgjdhSPFmJBxT5ENxp/p3fkDBb2P1+gc5ocJ
wel/8osrKbpKV5jjIQXUydKj2n6AAlqM1euZWMVAmMfL0inyyyTC1Y7fsoSZddXa
RSyt5vNNcvFPBHY0UhqeyZGcIy037I4iff5QTowviQA1fFqP+vkUBx0cSi8NVopI
0XpPYxjAnudYywN6dgFX1WSk1+B8cNY/cUqsmE94zZty/m7HuQKk38hEov5f/Xrh
Ffunq3XPT0IlVVv62sF1JobHI+xlXQpSf+JrQye5xc1YEnEGNAoBpLSvcL73rR+p
wNULWveTiNz87yVG2eT9tK3E2I3E8FeAVjobf+YrlJS99Tx9n0Y2TR7NEGSAPFG1
xRV6+IUAXyLpZlxJq4giF//I+12UuJCLHwjaIr0txAgRrQTwO0uXsbBgZNAwfY+L
RzJ6E1KSeynL7asljPd/uWER+oPMIcdMCYTHQ5oQnCtgaXRWuRUrGCSv7ie4AS9e
l/n7foaImCjlS1ZHMTtNfIAB+BJ/4njYNg/WmDaICWUCq1+nrjaZYGjo015XaL2G
3vW2OuYc05pX/sWS6dLQb8EbC2O0xnkYcBMy0zUplr8HJjheBBR/XIs2zPKxVgyo
/xEQScpg2BzYGihRoI1pqk0znwVKqp5JWm/stCsk1LPIxXWRi8q8jZF9urzXeO0R
omkdlZEbCCcdodkV+H7Umaw59pOKFrAqABNZ2rLVcuvLdKPBwYT/d/hOiJ/Ih7iK
vIDgEJNwp/qIdGpR6qCQb5Kl3786H0G92zk/LGSwW0gNTbKtlkcnzD5awrMs/8a/
/cmMRIru6SMNw5pZwKYErKkrdVQCNkTrN8Z+HNVphmgLp21FTACPY+ZULrWhS3JR
XuMFxoDKFy3y7C1M04doUuEjL0rRA+Ng68CCE+JULYFZ3ICF6Ge8WTHOkVlJ3+8I
BBZN2rEIQW20IrcgZ8ahFADKAI6+lyuXUHETa1Kh9xhWg5un1gVwT5VoPs4eKAXZ
UwjPS3Hg1t3fE2qwA2TPOTZ7ymj7P8snVdNRO6BBCw2ImBj/72rJftqXuCHyWVmk
rOx0Y+zRABiWxXacPyLIoVMjxNZf8mJlzclKonARygS5VHdURx+j3qfqLwExWj0g
HfuNFtGJ6W9WzM5uGuZ1ko1XfQQCmf0ZD5m21Fh6JEyyZNDySJk17d6/K5Ko7jWQ
wQH4CI7WN6WP/Jb7PkL0tPR0WoWZQeuIq+ZNdvLzO6p099/341JmCcD8r056eqsO
aR/Rj2xDvdD1vAZXrCF2GIT35atdkL8BhShJz+wXeo7Mabfs+4TkAJqIkVrH+onS
TrMlJ35gPoy+SOffBn7vPY3A1TY3/9+QJo48stD2vdy5CESOhCscG8pg1SBfJ9IL
o5el2Xxy/0wn8jb3iduDkPVrCX8+yigIWvA26AYiIVa42lEoTK3IrEdw8pMfIRem
jOUCaFbw50B6GCgCooCQ3YwF9tKix7Fpi6/o/sLuVn4gYS+1EiZzZm6enj3GrVl8
Pk7535Tn/23p769+oRZKeBuNET/oRITzbsnJp3qArGH9tPXFQuz79Xd8astzd/+y
oydZFW4fh8OQ97ZTgjd16sTG8nAcEOTmOrwgj+8t0tpzols58IVz4KFH7jdqEoTj
5pX3sT8Xzyga+M3EVte8lL2yvCFttGebRBdYVWiMCALlDYiCyQDLfx0Mb2wKJ5js
Jb2wBgjwUQsTp0M+XNMkOjhMn58cwf8YJ+5LivFf2Hh2arVyq0deoIS7SfnHUMQZ
PIWWllQ2ONdUoDjKlSOxWR7he6GPLUit4bpsy1TyHb+6r4bTySbkvzKxBOHT+hJO
nhMwEjp789SvPO1l6J6ns/ESYVbKWRDlnbI7Rcg84VSpbQZYPe2cboQX+qXUpe0O
CZ3lXq4+xBTsqNNoaRCUzR9BUhLx9I2iOAKynGeo1euex4kTlJjipnlzz85qqgMq
N6FpJ/70S6pVQpeR5ic+LD84Tk3Jb167zTp2jymVZU9W5cRfR+ZYOzwbB6xpbw67
yIsheEB9fvbqcrri3Gy/OFwM9ZTG1b98Y9wzi8BCoN3i3BYAMv8IXlgIBqmGT6J2
9pgRddJ9u/3JvpIvDGm9jAlX+T3dtkynuhMo8kXq+y17Vc7K4nbQFBkLigEv7xQv
tR+6DcGjv8fJ2/WcS1/Vdr043HGBXNHDGc1jkmg3wC0yr/87negvOdEZ4YBj6hSt
vqvc6CQfI8pkr/4oVXZYkpfpM2VTzEPAMXF3WcWb9rdP3k2r9+b6YplDxGcKygPm
pzpUsJHhy8PlY8geeoGaszfNwheVhKWT8ZZzW3kLfg7PDhAABejd2fu5nZWWU8qD
dI1LVzcI6YEuPoPLfdhOFMrF4NxvmaWDP9ZaC/OSmFuNsodxn0u25JoBvxXo05na
M/Bmk00o0V2XS1/kJje+ttZn989ip6lw9zc7x2XXy+WUG/Q8Yc/Wli8aJqy83Jq9
KnHxoCRBK7Bn/zV/6WL4D7jTlIS4NdDqQikS5Nu3LNPW9Xl6sOZ2ww/fZu1XD3QM
XsozIJv2k62SvbzcA0W8V7oUW/Ulzsu+hhf5r6dvKJZr83X8CE7dOeyzBPLILEj/
LW06ClGzCq7rOj2STXz4YypdXty7TgRXAfmq8qTcTQvCh2qyO0Fg1dcydVBG67KT
6xehM7gRzln7nAcB+ZexMM2/1fuLBhPYuDFcjqYNItkfDBm4uJD2OCB/SU8maIzy
zzByn7y+8Y1RdNlglgNDRsbaFrktzRjVZyNXkxfibOpZhNKTgR3HfgGMk4IGmEKn
Tf1j/vZmrcZ9qfcKSprMT7wUlofOcKb+j8Uqx3D7Q3e5GLrlQ2O9hnx9TJRSsiqz
T7X2Q70FuHmxQKXLPxtlczfnvxxRAI2M1q61dF/nhoJMvIKU60FYoQsdqfJnWDEv
Pckj332P/rL7OCc1zIjeEXPWNnohAhxhy2tbS9uUzExcG3u1V82/fD3pch6BEmqL
h6/EbCzt527/uV//7nwaJsMPxmZfx5TcONyLYM4tXFHDSoGbRYSHoQNqr90ckxOv
pFh7uiCWQb0+Uxzxpo9W8E4ppBRBlPZM63/2oRgwvl1mDSIe9uRh541MAQN9GAOD
cfw64hVZ4ch/xSltit2oPWHZ/zFEiEBv0ddOpDvSE3lpeHuZD9eAOvwhw4BMQ/fr
EfnXcaoDKo8wSOAibqN23d4WdeDqFPusbzYXG2WN44ZLt3n70yN91GFCQbobRnLJ
lnH+44Omqr72kWtNPldEepgj7vVBRgbUH0+nn0kaTQfLo4FK8qUERXPN+s55ANAb
Ghc6xqGNlXeFT0eQt9d21n40bKVw4n9XeHsjsABCPSBNxhrW97xHBbPz0bfE9xta
ECijiA4JSBcWK63CbCfq+KvcTtw77fRPAhRImZUBNZ+QmQR0i6dEkd9VLUAu75Ri
NBm4ACwSfuY4WDWn577I6tRkYqXOFbPhUhD5OmOyshTdY2beVRRlwBTP4MAVfsme
hwXQAw7ElGukytD9C50k3K9eFcR32nawMcDifIcwRbv1QaX3BDuztR6jFO9xxZLX
QpLqX7wH5m7GI41jwr6b3yRUaRkOhe4LvSxPGR1Hp2LZWmKccww7t5FSCBcVKNXG
nfZhfSOCbc3ynrf7k1ByT4gOBAgMjiQ0RK7Hqw9rhbeuILR5tgMGUDr5r835pTg1
8KWQ2BBtjitmyDqAfl2dKXEPcYhhQuMraFnTV7oqmRY0tjeA9s8pa3WOwALg+wiL
27FGPb/cCQi2ZDf87PQ+pgao2LB1bhPeWqrR8IwCrjWyuQzN/5FjfXfyQJqwBIZt
chRYT5YnaOZ2/cluRryXeyFhxjQ641mt0fQOkS7pNSnPTF9SSJZvzWg+VulKwoMp
u6Q5xbFNlRAxc0uDuWXP7M6QwiqKDE5E+IiyyHW/DybCXGnGBtKU849It0ONKzkD
rLmR3EcnacdLwvunPntkTRbUsYYlPxukKxDlC11UjjeIy/WAyUI2u8O8i3PUahuH
iKB3JN+hfs1GHSb5ppQ4j5bvMQFhsyr78qQhDkSkTuqK120g/uLJbzyBG6PaIMk1
fyeExudZ1LT34YYS9FEa8WQi7jwH6XSBBdd99LVmG8w9CZ63JWMTPbezg/XtLRmH
1Ih1XxI3MOoFPXgg2ILJrb6YB+n4GtNfW9NH51eU6U58K1uaaQMilQW2xC8/mUfw
DnbkQik3oKqG0O8h4PRBXKsouCCkIqMKuobSK1HyrkLpaHpPAMlNmczLCeh6XpEn
Qop6snruo3b5h1CLbLfxFBTe9amXMkio/E7JqnBI7q0fLCD1VkxcOVb6TVLW3wyd
3lzj8AGUEwujz1PQ4Iq2BaysMyLbJO/2SmMawuWDIRMVlvIUFXK5CMghJdlvXp5S
Cor8+cZkj4DrpNB8CLz8h9ChOVWiovm9WDZt6jStYdQ2rJPUWFzyfcPC5U4om1Pn
v3notf5CGQyWbJeR/WHHezM+CtQPxXtRFfqvEJRDvSjD5HuZK4VxdXLjMpnaBWmb
719fffkSh34N2UFXIrkJTDOKO2m3jwWXjHxNHLvL67gY3zePuAz03X2oT5E02hUE
ZX2/F8UMa4EN7V/DU96ia/icU3KIyhAywYC/YLXiFmImOskRJCXozKtztbl3jJ+D
8o5pOJvMumLnAk0ferAtjmnYUgF6LrNZYpPhZU0weayFVGZW/52ehn24uLTLZya0
V4oqJE9ofww4cP4UU/CiwTYQwIREh6wiC7DR+Bdu4bjRqshbocIbsSsRWBDKwqnB
+AcRrarkWcvn+BHaTsHz5/DFPVix8qhR9yF4Sdts8PNsWhrQfQ+PQfgfhP8QWDf/
0ixZYN4k/BLOcy8bGo+NmzuKngolI2Mc+RXU+52+2osrY7/RvtccKulLkyAYzLpo
CWJNIpm8IO/pcOoRee7BdvyPDQAYEGaWyUtyr2iQg3SC/YPnJ235Cur9NzksEKXn
/+prZRd3kBmmIWQ0DHaioWxP4zrkteO0cYSOPqpTPL7tsdOWcLkwYw9/wFZn0pEt
GifMoDxJ0JLPJb4gPi8Yok8KNF00AZsmA/fIEbosCeMA8CEoQcP7BR+Ohj6k9mc3
9c5+kryFXPYEDLdNJDzQvSLdcYSHE63sgVeEKoGmJfI9UbuCAdnDDtD6ffrcwAVj
RZyMZqZoRTnX4Rz8kGP3Q3Abj4DVp1H3nLzOLPr74k1X9wZ7yDG7y4/F1IIZ6shb
GF7K9bd7I34lz8wZ3GEl0rlvMHy1dqPlrhzQUggy+/xT1d0pBS5z6CRO3nLxjcso
bNFUEg4MWE8WN96hPFwSUY491DLb152Mio62DqiBhAtkuK4TzHHrU7itkFjM57Ha
OmptNaGTZ0F/jXxoefz9yCvHTypS3/+XvZ3YaSzTk6HUZ8tvZUSPXOqRV46rvVqr
PcQXsqrMNS+EyhUY6yowQ0qzURvqPYd1Z68YgXGZvok3MynGMiLcvHN7NxB5no6h
aEZRy3j7TENopVJAXlxOdQIHNcF4LfOWRIzUrG9UhqVhRuYC5hM+qG5aYTluucsA
upJPqky0HbebAWFCDdH201nsh9Z444/oC+H7XobbzFf4EMa4YRKqYPwR8zqaTVl8
/9+OpDHWr+Z+tMJh7XJM5dnp+I68ixqe6yQ4oA+mjpJlydCfXsODZdl9WjQoIu4v
qT3rDWHWJg2BhX1wiMwyTrbhbb0hw0j1TEqP66s65S3PZvXfFxJh7g9/QN2Mi+Sx
N/B79W1iH2+QbMv9JpQYUz+LUuZeeRDWqM0GLyU/grAkAsu2+70RP0f/kfPgsIdb
FnvbUmQnrRhMJtin6Ive03qKlMcIaisIECkI+Ic2aIMJYm+MIrZmzsaMeS1X6fvS
VySVXKNpmCYC6a9DyBj/L7pZSrm/GrYsytSqfQRgiqDEpUCwFbLHn2rFQ23/4cI9
1+YNvpnWFY60VyuSt50SGUxaUqykTJfxP4zFJfcbrmjz4U0I+CR2RLCOHFY+/HBD
N+4KdZUHz7sO9bgT6sMmK/YnsqIS+exM+4r+pTCqkt0UXfIGtMuSpfEYp3Gzso7c
j7p1HlqaWC7BYPWRB1Wszy/8GePaJR5XhjI5qN28klkvLvjfhvO/CP9ZWv0KfQYw
By/PBd0lhi++ieq5wtDD5T833p/DzvVusBzAINTY+kWSnnlLujLZcIu8Cl3wK9GG
R18xPS5T9jIYKv8e1mVKCxZ7botc/MHVHKtaGf3Ynk85E+TdR2wPEOiXvtvR+wI/
QuR59B4jYMEDNNJnABiZjanbdwyFrUI0hqEWSW6571duVZ2/gEVWh3bMSkzyZpiu
Q4SXXP/sjTymxuvFjISZjqAqnwyqcejolwHj120T8lGryQ/b4FEl1S9iDRj0Rmta
eclB9Y+tDCwTP1UtyUCuK6TYCotWFgSBDDU+I1pV5Wigh/+o90awhjBp/CbiDwEt
HqXS2jAf1Pvfp9cCJmMsLpB3GA7gLmDyiAsXEvSavlnEJ6OhueuCtNULwxoz29qI
aBC0rSv0zzXkPWefeUZTIwL7KESw1tVlEp+S2ieWIkUs2N8k3GSWd6byF4AwGEG3
K/2BzyWyIiKBiJZZHRz8/sNGDIBF8uiRjs4/r3ZRa1w/DFJuZu8VbM0TLEVf89GP
kkbuQ/t1IRJKfVpHn/tloASA7lPDhooqPT4+49kRxNqrcciZwjq6k9jkpg+guLKq
1NBT3atDL+mUP17FMcBiVQm1BzSEW5UgD1cahzKU6VdSz8dN1bUngRXK+l7xfn7k
HIBlJemcEF6QQ3T7AfN8VX8hC6fRJ2ribFM/ZTAbdz6x/Bt1aNaVIKwLI1J1nG16
1i3rD73RAFwLT6ddGiEvSSls/wtvDKcN8DolE2MnUwaviVOJQZu9vayrCSF97snB
hFZhJ9EGCirggZCPAEO7FMJq3YVf8WsLcsG0xLUjZr//pI6MHRAQLMAHBfIMkCH9
ebADBZE7GoGUPQbCjU0xrQsjQMewh7E1ez9fV/HqCxVfKxVUXuCeSKaeIhSlj65l
V3B17qKIh5HFuoaxfVj6AcSgRu/p5neVhy8IUFgryhtxwauW7Zv1z2Eoijce814j
laNDA0EuEq4KXTHQBOKzg7EutyuTivMp+8TmGhK3N+kuJU+Vsh8VaFzHAAdr983H
4eE3QBG9h3/esfY9fem9gVRiMj2DPNmY2U1Is136hqJ0N/M5+yfg3VxK5F2dXx5H
s9ZEnHpUcSK9W6BVGw3cEArW8rUMNFQ+2rO/YfsbVTKUQpjtNIJnSY3k8K3qeBfi
xj3adM/E97/zdHdReXxcV7uK/3c7+D1aKtb0Xwcfh6jpHZBzPpMPPJOSgwbjVfFv
f4HUr9uI5R+f6LvedlL2bIaB1soi+EsdSc6Xck3goeLxiq86TuZGAfBf5u76ETEf
HXjVwg+xod4ZYZ4Bs/FOiu6bwS/lCgkG99iNJswGKu+8zorzT0Vbnb6Qs2Y/4NYS
x3WAcgBmkcwW2bi7V6QAHnQcoC6ams3Km42WbUdIYFDi+aip8da+aNks4OWDbKHB
anA5m4MA5XV7uugdgoWxQc2czKIR7cc0N5cKI0AMtQhjqUZP6nI23vCIOrcRnNcl
tYkl4KlwJIw6lbcXVTuRoXwene6KKFD7++LbRjJdzGPtI8G6Y0So8av1DPqPKnm2
tXJRwVsYBgDipj6hQ2vwzz121k6kKeLuCWm2cSY7zpRYHk6duk2GT/g3/Z9wTgRN
/eC5uVb0kdCUybupeyRU7lQl+NlmKBc4CrgzCxJWkUcSpl2pb6QyQVph0dYEwX1h
vuFdzFJKWmLaZHZreBmN+2CkTtVaAIyPc/qsso1KwbfYqNAIzgUhguKuCug4n+3z
W2oXhTEJbkNyc0KlBl/SKn1b9BOzjCN5fYUneu6H5Ea2ahH7ND7hI8Tn9r4KxA4H
2qnkh8CGe/xW2KuqzGhdJpftVkBYYm1l6tG5E9kNA8mlDpg45fFlfGwYcUOy0gqC
8tt22J64Ef0H71odkz6i/htf6qut0tX9XdY97SnSmVvI7NtxMGtQuKozj+41MEJV
FLXGFGf9JZaBQ1oDVR42s+C3JwdzlI6lO64CYMZp5D7h/75oAjb466Q0JZCdiDgX
o1uFZx08s/rKxaoomuWw9oE927vb9xUGStRfdjAj7KdG09dKPbMhpJRssDi+wltD
yhfU1Ph72geioUZ1ACs2UM9BWQbNkPMiMzdmY+84Ku0dRy0CkTaN2cV6PVIYHHPT
ORdcDABLpC9paJsQBRnJD/3vPPIC1vFx1j157O6Gcqlr5rGWkWsm4cRGfoSLpnQn
8VLPBLgK5imE63onzQTS/mURDCYdcmWNRpy+ZPOyefiOwvGCwCzvek3wN/ERSfOF
xPU1Vrxl4QWDwH93NQ88+Wz2p4waSwiLcXsBYXq6U5ggPLo6Swols4cgA4OmeSrg
QNQY6GFn5OkmqmGKJmCxzE6/PQXDjA5bzZ08jIvCS7Hf26hVkFE9l63b5lxkhxog
JrtSvOrZBgPEP28IPsBG5EkA5uRV9uPokRuPsm2neTTvuj3TIczs6XnleJIsaYAv
dF75DxGN+Az3MJjNemgDIpNJ4rEvwJRWUiTxBG4XzYlXvLUaDd1IzGgtMNa01E2T
AgAGqgLbN4yJR9NddsiPWbQsm7RTLYZnHBeKPYEDw/8PdKz8HrD/wFb1QbpR4dJt
3ueTTxaF8LOtv7REzqVv8O5xLRaxIoSn/xx/QvUJY2edzePUFLKdsG1p43g6hjJ+
PJbHxxb6ZBai2mecveSu9N0FpRU7Ps7u4qwPvKexg8q/AJMQrhSCWqUOPUbTYzW9
allWrz5kbpqlX0MQYhcWNhnMztWBoF1un3PdxI1mCDevorMrzoi0xM2uPXMegFeR
QUjdaBlbqhiuEdqlVGYxbIQt8qTHxGSUZv8cMToyIJw5SrRbBCdncHKwuVb2Bzsa
QoSOc85KPRRGJmvozY+4jPhIiPgvV+Rume25oNkBDAYjXYXVEy1ttNI45dCSijP0
H9lzYtT7B0z6V9IZzviPs23OW1cqDbmTE5/VAZAXfLKD8DRuIfzP/KxmrS2nx9Sv
hPbtf0YaEKqUkGicKXpfzJtVx2q97Of0wS/i7ErURdVV/sTzg5FZE01qH8Xe6F5n
o84zSmYM/P177iqXakndkcscrv+WSM7/3Csqt0AvtKkXQTfdT0GI47j1WZiAOeys
dAxtxsyvY/FbrwpHpJ2LuD4mK4Kj7+Mm+NBOWrhuH8AfaY3F3eSUERI6i/1hSjiq
rDC6fxLHeTPLbdccmiKt29xTbKaQje12PcbBzWtvpT0f02a0IcoLy0eAuu4fihKm
jCtfqa1uAbSV7LQm87i43L20l3O+aIeDCdTfLmpoYLzKPKlQhRZcXve/MVD0xRne
vSeCS/ms8aXAjPz8MgdIjHwOO843hjUT5bo4QkOj6oee4w+tkDVHmzwmP8ZZWhqS
z3z6AB05SQan5DQCOTEaC05BnRgOd7Tw22mUavVJvdd7vlCN3nKXR6zriR4gTtRO
E8waCI4hk2L+rDCOwrx5xyMtpwBhX47M6WJz8ZbWPcpJqNPp+8stHy123wiwjoo5
/cCqpNfYTuaYHdwKcq0XbDqA6KqEQqlxcDajShSf6rJo2nqZ+k5ei7tLcyLZpp0B
lg5RSLhx5H5yBoeNjRUmfUqg/ndKUwiUb1HeWGstDk5MqkVv3M4yNLaecm+XDIU3
g7F6huglGAsePBgLfZJpfZ/k+OGuY5geDsH6vXszmKl2EdQU7BHfrFONj+ClDGBS
9xz25e4i6Zxo9IAJi45SNnoFq1qNQVLWnJ6SMaAKj0UA0GUHQz9vKY/8xrw38RtS
Y+bvP+cvF29PE8yiQj0TCrVJY8IzleVISBnDjqPXljfKXdkma4q4QEeeHBT1MQXs
gsaNAl0y+RfpX+9wQI1Z9xr5w8iKzeS9/lttFe5yxUO83YrbpE7CrKcCEHLcCZYx
giinzboHeDxyjQ52RRa/COS/a11huKY6gl08l37mURvp9fdKbYAxVUh9PgGKVBxF
B2bc+a9o8kheRAq/rl+JJSwa18fj+zxKj5wubkBCx2FD0OleyNZoqXVgtPowKu5D
gi4nYNm8jzU772CP9ljEC29rZpHzGeaZJwIymgoUTbn9oLmb7bV8MfJM5fHyABt5
YQFFyFiYv3Jr09DGObxM5ciCF0ZKNXoC58gGEu5bZ05unSs2ClPLE7C5UbhCa/uS
eI517heZ1wLYThqhBfuqogi6TuG62hyCBLHJ7aPnD74V9XHYX6aHVD3raF80xlGF
15gPIuBcnQGlwdjruKqL5/8pIHwzqRTUaX+Ai/u4+QBdFwBazLNej5mgDl4HYsSn
GiT4c6kEvqdyEfJdu6gFUOFDRP82ZLQ9bxmcFleyiSi89j07cxQdgWu6G+8pyPls
TapqFvrkTxdhUxIdNZKE/w+uDfUoJ/PtWFT6OVnsqR/sBZbl0OZA9pCEl3838dNq
7YDGrNEa5mQWmxpNzTMiHT0QaZCuiS2uxmnEPd4cPYep74cWcfQBNTiezxCPE73o
MG5EjOQ5WxH3NlAtSkuyU/2T8sRWDwAQcrfqn7hOk5uLSvH4moDHL7/xRjWeguuQ
eDHk6lyZC8Dkz8m/YONAI27JZF/er0EPeKXkXK3jaDkjevXP2ni39KnjOMRfZn4g
4VQzJ2HaHpNGo9TA3uAtYuVm8eZkQhz/p1snwACVXqaoW1J8FjYqMtg4YRsO2/LD
KrCAkTIWHiHKTzbyzsDCbQr8V9eCDkqUT5lyGhtjGodQnpPMFRvkuhYM+8pM19mq
O91nFQJm9WdcInnGBd9k+oHTq8ZpBjmLBXB0XITiGz9o621HlfrISvgzfJ1tSbWq
xnkdIEGbsRPoEbKX41nYoDlcS+1jXobgZlDGaZ2iaRLA4EgVCWs/rC3LTrUtXO07
K+F0D4Eak0ZK5lk5rKPLlZnSSpOLfeh367y2iILwi081V/Sd7bg0vEHt3U/g9Ber
lJrnNPUkXalmLFU3qNFipHglLZGdSaDChoiF/QwUDhBh5PkoR6oAYsjdvzA5/Og0
boGDcZUyOynD5t++EJyNKQNBVuSaM5xsnjhT8ej3DAH2/YIaVohA2N+4GXrylalw
P10bKWyG1epJ8UMS4sSrR6lo1BVEt62rN5zxhwKawZoT+qb5cYXFVeZ7I+zBW4o9
bLHn5aS6BPdXCYeAIEecu4rNbi5UybzpD5xVN2TxF2HHWHCzWM5kkKUe9QdynmC4
PTGwy0OUh+Gfx+9qgc2WFQVJAhPy+YZ2flC5NM573LUb8RpPuQkjbnn4WBETbOd/
e8d4QklTlaTJATQOTm9yxes+XUEY2DkAvDz9oVPy47o90hCZumbjilSdNDcf7g3I
iU/SV5e4/Dgr7TaQXHoHQh3wiUvXA1BMbqxVvyVvFhhCvyUw57HoWJldvTmpr+TR
NmReI8Z9Bmp3FunRWKlToXtPgZsDtq61MPttbseB/lFIPcFWd/DXO+8xL2i2qNP7
nQMFjIURlqKh6NTLjicE+2JH2LiJMz8R7dPL0zEZhD1AGsfwD2kXL9e9CzxNtmbM
6SAdRMH4dlFvGd3yDVv9UZUn7TD0DcFHYQBX1pxf25Tq+7eT+vr+LD17iGDq+qVG
wzj7W94iZgzkPsTgddhi7w+mzcTvCWGk7nZeaqq0KgJD/S+MCZg/0TW14501ua3+
EXDnmA/TfVWhhiqag+/arK7FC+sHcGcoWJzI59uXKF7jJbtCGAboWN9f7MhTJxl5
iP+x4ipGXkpcfvngu8Okrz6vJM0i7AO6wV8p9BuFPTt6K02ZS8Q71rhFiOyD1LW6
Uar4H9kIQv9NYq+YEc2lGvUBQ3C5/YQy4StoAQUGICc1gUbI+9uK12ygNY1RH2gw
E/I7DdKZYrxJh6MhS+QISW+lS49CeLfF2hTwu9vcWBDnnYqmCU7NE3/DkAn0qLI6
qZyLu6mxBV/9VmETY8i8MihGrMEfu85amL14O+y5Hd0t5aq5R9DJUxBpEiZBc+wG
HA540C3lX2eFfgby0vcl/U83WdiR7G1tij4KJ4c4YWOxCAwGU5gKgLiM2KKTdV8h
ac7SJ8kQJQczYctdITNFtBDz+3rCN7F8o4q+ghQQVX6uRwYWS5in5Gku45iOQokr
OMKpziPqnMBxOCrB31bB4gUpG/ktzciICsMnq2iVox3XApRM6exPkCWno/t50+Yf
y1jiWwG7GXY2AZqi2flV90mRTGx1t6QBf/zUwTN9+1/9ej0N+UWwFU6ZInTN3vGE
K6FEv39OoJY0D2W4yDfihnweSjMOioGaBTSwdKh9Zz3a7a6q0z6krbQGzv9Y2jL2
5JJl3EJ/R7pMQ42LevPjtIe79wz48OG2+/ZSxYlCF4aCL/VIHLOBqVMU9clCSMdn
fM+OpWhs4tRx1EoLmip5ZB7yVOXSrFgr+gpaQc1Zuzk3y3TRoqUwgLGnfpjL2HeB
S8hWP6ZpocZrj+/WF3wWXwqY/RnPvSU7YTvdbzNdP5P4kYdsFTIIldwjcPnp0u2z
NEW2K3YXDWILYU4XUa0lJg8XBn+I8FsmK3LApzapsk1PAkwfQFJ5hCz7GXcQDy8V
aEwYNcwnBfLcveULSNEKAuIsogHwJbsxxea/Ue2D2L3KBjeuNkE4foUgJaIMAxc1
eHctsTlGZ3Q/hinUshG6fU+9/uk1Q6nX3iEO54tbeQI54o2sB2aUS5E5IV0MKo2B
Hp7ina5DyFWPtdxx5/Y2qP/BvlEVThItFEf526mtEyUKAob7363zI8YUGDH2ilvX
WHnZtcVRbr9S52SmCsYRDdsUgmC82jM1KpcA0q0899DKkJvKIWcb3NiJrqbb+fUL
dO2XX5FPeFgBkt4VWRFLXeWxrUItzZL8h5SiBMAfKlmnt7k9eRZTmGmFvMhOoet9
aAEvUUGQkMOFB+PXiB9VbnM+/jFppZ+Yd3vLZVj5Il/IxNI+qSPlAUzKgZg5uZvB
7E3TOekBrq/YG4379r0bNJAn+ezejGboLlFseO0/nnzKHrzGJc6rJKGAVzbhyK1V
xNNLpAJf7H52unSQL/Bz30HaarORQmdBI1ZtnDTYCoCqgIwlab+SihawaavY7M6r
/LUUtGEMcdiZoIhDmjKMZI58IyGO70W8qmngLRrN8q6MC/OfbD8ZnM74jG0R/H/m
eTAO4CMoFmHC6ZJUnihvbHFLGbe4MgoxdVt9eEeZnGqRlOGDklwl0rAblmd065Kb
kANcBhvZPpbe5maYd28vK99AIEUT7Am/sY72PHsw6EzT3hrRzNBeyD4NHRPB0/3e
E2EfIa5LdAh5RTZy2VtNbJgGLNAm4L+GDV5l5Xv3KunMfWiiaHQ51pOeK3G2YMI5
bmjDGtJDDuuZRo0nPgbTj2F/GmjJB1IMil3Gq8exb7F/wfPEEgFtiSrizdb249II
8aaPRgX+to3O51TbQ1z3ys8Aj9TryDlDreCT6ftLC8c8aEpm6HdNHcJjNDV8LVet
ctCPY+knpk9I1Q40xGI5YjExjteqGx8zvxOmVXbMNctymbEXDZcIZpVRiCCLm3lz
dJW9jyA5jlbgbNVSbvdTuxBO+SGhvBuaO2pCM+B5ZfpU3nLhltDTh3xwZjQh5o3z
rxGY4TW1BkiTKWB2R3+yy4jTQMevZYN+aHihUstir5nZyLrCI2jZJCdd0BM2EXoV
IJTKfBEAHwHeBABrzR1cs+yNS1VvQ8cfMZi5x74jaASEmGXXdzJgQxxMOkIznB47
Tn7T/7eKloJsa+EZG3Q2iZ5SBcT9rC0HSVL4I2r2NsTIaXtU2gwygQuu/a3zz9cv
cvpOJeIAEsL0bl9OQCxxS14SjMEnbaDmAF7FZta2jpHuq8OzU5aXNEk5m7fiwXhK
Uue9/9zH8dABdMqRCIFtz6BQTojXnO4aX30fbhxLV0W263TtiudIpoPyYXd114+W
x3J+QggwoZQ5vn97oGl4e1m7xZboe40+pcjTZOGsddrnL3RKRT9285dS4ctgxc7m
E4leM2qQD5cMEBFpp+ApD86/G8kugsqgKja2xaeufXxkBvcmpzl++7WC+4m3gU0O
Z4/QPzYYrgZVdtxONo2K4VIve4X84XQm5Cy1BFetLLbd3VzE2qwSK5XGi3258w9j
3mtnUVFhZW0LldfmBqEiFwnI3T4Z0Fln2MEEExJ+OoCuI45rQl4KxD3vtN2d/Tr5
tRrIMvCkn6uynB53hEFs5Lqyp2LzGLdfpDTNAoIuqCsFaQKnKsxSkV7xTqOr/S3Y
nf4G2MTEoxlUotO2tUxLnOaE1+X1OqbwZFR8Hz8CSOnAi/3mt1RBTFaJB4txwchy
LEBzgwfJltGYb8PYRKwHyPJBhNLb44HhKB0hqVQYSJbhciv5DD/Y0onu3Mg38m0w
dSOesuQyjyLmeZpcaNtLdClAbath8QI2tO4/TbLwp3BnTTXkOwFQUfGdN4t3su+R
IbM5yLIPueB2fWOJMpVDvfKIX3Fl48k23F9gk/pOcpHKHm+Tt37F8J8nso6yPvpA
o0FJi6bgP6giKTnISrNOG0X+dOqTjjnhx1t5SkkXXrBOFUzRPlqXIzIwvvjhotq6
NaUVyo292LhaxX0VE95e5qUOKzP2uGHbpYappgPWfuI9vJR1eDUWOV+6ATMNYzKs
PtQy25efNqJgnDB1BSCT8FzsQKDy0UCAF6tTT3Dup8iCk9310Fpup2+Mqb7g/KF4
qsS23gH9TOdcnEuSaq7qNQ8De8vz0GZaJP+sx/k0iFblxdKSILYhU2rGC0FDrVAm
Xjf6X+Hw63nsUqcql6CWkEWNgdLsps1Y6WrHpkULq2p1i4+T9rV41A3ZOkG+I4Vr
u937ziYFOxM8q0lo0PuQgU3CTBV9UlQ4DQTofa8+T0Mhp4crisuU9m4UbDl0T9hz
+1PkSCT9HedvfcVBXrCzTuNCDiBgtE2bOkNn2b4F5qOUOpqqubHqFuhktPCMZNIb
B3KUmPaitOigKL9qD/TjY/LXjT43tLbVLR/xpz59q8yz8Pq0d7VnZzLlewtk7KhQ
Jwrt+TFvvaD0ceqpW6WBTNWV+DAyptvZoAIxzsro8oIcOm9Z0F9TgqxN3SvpLI+C
OCcMwLrN4dVydnNx25oeJZnN9Rb+ZAsIHZ81ENzz5yU1EaXk4dmi6QSrBPnZoxoM
nsWPo9URX0F79khWcDXKr/3yW4EbPAbSgPz4XraWNcnJiQgA+idukeyH1VBwczEL
tuYBBm6e7+HbQHbTV7yHESg+LuCxiHPZdetBxG3O90eci899Lk2Cvt126A3n+rI1
vic5KlRrP3o1crHlwbcMG2112bV/1A1b2TtYezP7NdBuWHuSOk7PLgo1xJOJvF+x
M5csJWDAbloY+3ZN078TBnnVtarMoPfrMOhlkUErAuM3Xz+hO3oLDrrwRIG9U66f
aXvB3TnEdE9zE1q7c/IL0bI1jGNmt2flPV50iH1r5uw2kZ+b1K/aMjSLfI7BPzx4
1aQ9uIUD/LF+HRs+8XtWeYdIVr1kC1Wl6A+hBpIEbwQO5371Z1MTT1m+uzXWg3kJ
zJD/jCmXlKNpdM58/o16JCYixodwVG0lPLLDY3M9f8lB+nMzLXspUalLuFc1ZFQy
htmyJ1ieFJFLwefQK+D14M7r7K+z7PtWIJrTuHMg0yh3zHmACGc7NAn60rHtYyDD
/jfJuR+tDd/1mVwuUlnfzOPERTLm9tWJn4EeWt7qX9Rtltaoifxsy8dNfEKcpmvg
91uv8CzipTG7XCYBL4TtUeKAX6Beh+EwGVyh97kB6JEn4TIgRMAgLwO4NaW+f97u
5DLLMacVlda2HmT/ASIilaluYGwSa/QPQwgWKSn5ddZqH2aLtb2lmZ30+XCBMzuq
FLMl/spggqpE/v3SgN0nhM6os8zvTyQ3mkM8fnRH0fAbiTYHLA1dL+FgWZL+1pGR
zkVndEAnIyHZNmJGZBfuzaipRW0RtPVzjHQgpWf18uivyXn/kkX8hNQHomQxY6F9
liEU69mz3ZVHUkNpGOSHglfqJpwPP5paO/brEiLXYXPUNd/WOzoQeJtRH7u6dLPo
0t2qgpVZWQm3l349lp0iRfD4mSIOEooo758d7kToqVqhM0A816F/Bm6FoUQsMn7a
RvsUI6UB0azzS2l05FslO+wHiNdiG9ArwVsaxFQLVdgcSwkcos2pkVcCqFjrhD9j
7KqGNSaGt/iKQZqsYtsxCV6ECvG3ie+p001gsWJYW73556f+4KfxfeUORyUMjh/c
PcRkMtp5PlNHd1zJHHrulwVSVMy3W3ghtVRVvqyR0pvPBa3vAxtdekEFrw08vzk9
oK5qECxGyoU/QDx+B4viD9tHbrlHqiUJaGpM16E/uKJlgehk+wG7nERxyyf6Orjy
f3GHDEeVMHF8z2kSijxStXhbZOkyiid43M6nZa8dm4S76VWqNAErjFgb1VIu6AV/
Qon4+06iqGAhDErVOprtlWFWsB8eiUlXSj3FQRhYSiAiYGupABqSwTvWq/wQ9EcQ
1wKA1eWlWXh3W58s7PMyFIifQFDQpk2Kmu1BnisO6iXiHNspknH19l49zHzOSexG
XuEfOpz1425y588vAd5+oFJ1mSOtbU/kVZqsKGDp9rR/pAqOKgOI/Cozs8O7Tf3P
IsaKEeW9V27xGs5r/OfDd/xpP9sanELzc+4v6/ZtPWz0QfR5ialrfjX8lHlaFj6p
vXzSvT1GlMecTkKtfCReLAJMa6ZWc3IqGmw3GZNAAq4gx4iEJQIzhzzvVxN/4MsQ
V97sD2ixaoqJNgsx7W80XimMwoeMJrsMp9FVR0oaiZF4l+0P9xZ4rajfOzORadnR
UsDrI8bUrcX+Dq6bXhAcXc0f06HDhPPJUkby4208LfDjousA8l8WBTyE5ZrA07eI
brBHp7ASzvTGwYJqkqW9h6IbymQ7A9SJ2ewjha1x5GLrrlKfWNIS5QNp3lTRrdJM
n/pVij55sX7IyUlsR7ItY7bFh/Cef7gogJ/je89ezMU4gUlUOO3z9SxlvCFbkupl
uohOC0dbqLM7QZxz6JezCtg6aFGpIncaZlUuwxWSR8tMiBR92HfjEEieFekauZgI
Vov3S2Pas6vYnR94GqYuj71Czqh7StiivnF71xUQJwO1p3KwotCA4MYWBrPpPfiR
mW41UtEGJhbJLd6V2Mgomw4v+sR6ws/GEP+tyQJltP5ihnq0kc5LkjK/bTkF+1Aj
h27Vu40/F4Wr5V1glFf8vrn887STErZjaZ13BAefM3p5QcjTSFIHNoA0ock+ljWW
zkSBnzv84bboA8lkACadBk0dxaLYsX+VKzVpnJX/wi3o4FYnt65KV8/5K9GsQ1ji
20dblKOF8U7ODiC0ejfQVOJSKtkPY1FkNcZMWNEPebLa8wPlQGXlPH8hFMPIhyrw
of3lqLcdv5J3bTDO+4BT4uLX028udQMZsGTL4ZG1NtJqNCCSvAikT7msbr+eFXLC
5+ruRBLyZELixBPAJC7KkvYiuRorPnLJQ8KvdqIFi9+nqxC4QEWJfzCLZ093ThN1
yKrZuZa7k0Ccmz+y/hODuyKjhA1Fjib+xpKh6Ku8ldy+dMzjleH4CO6j9OqtJzoz
vTdYymXKHMDrCsj1AXPBUizOk7rL424Dow24BEcFP4jf8EgjrlXcscWu7u/o64Lw
gUfhC8hzFMroNdNIV0kuB13Ol9EpD7r+0x9fEgz6M3Dzxdg7BtEqLEy0l7Tr+Vju
LdNu1jwK3tntGJMjIV/hD4J+nf/IewOau7/Qrvbqi+WW+EdiGb6zFEji6CJpAbef
bPo2vRBlEiah1dqHHKWYI2ZvAXWor8AdgTTaQycrxAanIYPacfRN5T/pKEjzmKCM
3brotTw9/7rvaToCEfIr5oyPGQhDGU/kq1I6Jxy9J9tTkaZo8Go6TWycYzT08MY/
Y9OAxUEWynfuBTzcuZubP9GpFpcfVh31q9npTg/CIi6paQBVzzfSMIe+o8lyJ8oM
kzKjcN4AP71Qf6jYk3xOFG2A697Py5dv8x7hhN43ZJa49HYZlEpAfCLUsDPzkO1o
ET+d1zp/4Utz38w/FyvlToeMypE1bs8jHxQMfHJAfyvri1exJ4y/EqZeChhz8Zy7
jSKau2kU8s4eP7ruJI3jV07JeIwx1g+Q7RVxSi+AHt1Ht0nePptMgctWXb4fflz3
KqfuHUG7F1VvCsOJd7Ajnc9pPrzR/+YMlpMAfpRlTr354N6FPSNbCgtbejnbFR3k
boVu1gQ6DFSp9gPe89aeADVexCldlIKWY9srKOpJmECElZo23ze8BbLTRyK3XNTQ
0Bjo7PG4SEPjMrHPJY2qrgB1XtZk5wy7dBmO9Duu4FlJOKuTj3gvBDwxqg0c6CWE
9Ojz5K+a17E+vwY/sd5G0k+gAOldirWcEDygY7gkZW+eoIjOEKyeliWCYguOyRIn
yNRb8ppSmeqtfd4hi0SfJ9fe2Sa0s9kjyvsft88CSDy3HcUoKqeYivpnvcU3b7CW
M0z3DXFfag3HYzbIJpoJKNzjX0vPAo0BWNT9ozUbkg0W9TWnawNLGBNk8M+htUO9
a7+AV7Gdt3KLO1/BugcRArT3QzDElDMB6UdJ2HvwT9V3R2hTV9sK/IER3dzL3NmL
yCmO074f6LV46IlWfdquOSQbREkorC4KlsmlNE90J06PvCS/J71DB8wRrE6t6OMn
M/lC9NxXwGxjq8UJ0++cun9WueziDtJ9tatar0Mksm7mryzERmAtq/JmMtMGEtep
nAgAA8WQ1cG+3mJji3u6VxvpYz+eHoJ+Ium2O/nzaV+5CnoEDBoAhISelmwz10E/
PO9o6N1niyZFavH7V59AUk+2ZJNxJSAbsffd2IHZ9PLcHfBc3jNYwTxaH9L9mwpW
7w+KnMVY03b1MGisujYssonHbolJLZUSGvMDkb7H4uPnq4E5Gtpp796J4tohVUmu
tKGImqwJ4VJjd/LhIkon9Ork3ECfx0fCEgWYSWTLKObK+7uWLIdTNmwMx2YK0xhP
hcQTqNoy3HEf5ACqF3gvWSD3H35VjUzBqaLmdzVSfiXh5gMiX18UjlzJWm5TJfba
f9RhJgjUfRHOEgJDB756erbeE41LG4rLzXadaI7MN8NipFuRbz+UH43lTsIg4R5K
qhMFQGNOD0ZlsXM3Pp/kfLWSekSxQx4P5+ZGAGumT4GtjUe1oCeJL4GmTsTnm6aK
8HvwQd0gZ/6zHyzgYqMFA1FwA/xKZK7RrSR345FkswJBcUuibB1s17xKCNTza1DB
tOVLQNkLDo/KaXJMp8u3Ttg4+PkUM4ahtYFCn7PYewzYBlHn8aQ4uFJjlac1MIP6
Z8ibb3QobdpotyMq6lcyVKU48OFfUwIsxnxiSUneSsxWE2qaEC89jrWWONgYYyZd
fQoueQ6OaJW+Zrnf90YDMR/9cmclUZC77lCqmb9Bc31OeS8mmBWUDls9x4Prsitg
13ZdkPoQ+JWEOcM+Byb670YBOuYzRikpIrkEvcvAwVX4FxKJdeUX2CPBhkdXR3ce
HYiVaim/wjZcXPt4X4yrC5R8dqsyg7Je9An+2OJR+sSDbF6w+8+v0OcdOf0fFjSO
DXe5fF7HYbks5DG104p459815xSRAOFh+SKWHIDAsZ37WwohPjlPQ3vuYcHIj3Yj
uqZo6PPiNzGi9cvLBS1rQwpKhzhvVA9dl6oNH41nzdgTSkxgM1PTTDpYQDDxpp8Y
YFLbb/dE8uB6j+cA9qIxoWgtH+cbuEUmEU7FV/ZJ3j7YYbM6RJTL+N9fITb+03UM
r0stCbZn0Lo+FlcEmyQfn9NqsOYmwqIUHbvOU20wsDJ4BP7K0b5oBLeUkrsZ7Qgk
cvkdUVVqyPP9LG05ba20f84DhQBlXrx+9Ki8JIGebFUSv+zSQczzXgkEeyzVTjoz
CLzXY0mlm45hQ+5XwcdufEwZMDGmNTbV8xLWt4y75GXVnYWUdOT3mX65LB6xDbCP
obQ0DlGSx2ANUZYcT/4QGAY3PnjZR9KuLd71swSs/4h3ZD+VbWB7/IKE+gSMaTmM
N/3+TmhD/4l8u6+U0mZuxanW4oXick5Y7czvT1yujN0MfumxtDa40/L2IX+T0w6s
97uZHiSFMpjuf4c52QbMJejQ7B997VETiUlepIQerYDFZsVgtlAhOVTXzUts9Za4
j+CWc9VpBs9XBbPI4grejOL+SXzTXbJ4DXoJNdBkVcB9sI8zuihnPz8oLWCKKxML
RNpLgDdb1iW7BH1EERK4RjoHb30mRKb2lrDrcqSoKeGyviQElOsmchOW+Zoob0CS
0pZYib8C4fRUu6vPJPqpIegoi6Uhva8FpbitdCaP3M2Eg4fwiYftjmrOTdzf6yTl
yRDkZIJDY91uhMfUlnCNUg4koPDvT6hGnFOfOel3+yLJcIbdjnTc2QqfXsErGgfk
06xfBvHmwbyS8l5B637rntuzK5gtzwlgsX71SUJIuNi9Jn0zW4F/UhQJUHya0x1X
MK754TLJY02VAtLVlFDyfEG+FbuZT9O9qiuhZwdOqEcqjGB5UwL0sHevgfOHGtOr
zPm4mcvAKDVYSKoy6KZgo+jTE9W2LZc/8z6N4UQWDMh+esbfjTBQDKGXYy01spY0
hjWFDN1rOHd4V6442uURvGfSsZZbIv8p9mxGmk4zRhSbS8ISdMBB9w2Ug6+3ecD4
jc+GgEiTpG5p7E9iStbN99KDpMZyNfmMx9DXiEjFOlIJ19uWR/E31/TUXdqGMMz6
99ydjVYE6pCBPSe8Ac1XHAeNEuXf6YDImjBJZ0io8n11XgGMtCCG9R3Zu9x9MRtY
54zJr/zHDXbMVHRmh94KSuZs76Dn9HuQJoVMnDUJms8o+gm7J/Q3U3uubtL5df4m
JX1XOtaCQulramXm6xv/ZqrTg6dLsWeC2b7o65eNPfqQ941CYHOt4Hk/NC7Rti3G
8+lRigYax4mB6HBD7hJTeKps0yz4MMNd//5XzdD68HMn5Y6zsGP7APPXRJ1/dN+n
6b10dzqzcW0RJR4TNS+of5PRs7J44G/K+aQqRQcmMMd1Rl1Z8z3mL8z0Rc/RHr57
YlNLgRVHal22O7Sm1ujdqklI+KRFLz4uxfNZ0k3xLcKDfMDxs2/AN0Nz98QqEPUB
iPyuexUFZPuYvLDFHYykt27A15uyzWWQWC2CKemY7aBs11S/TRdPHVw+oPASCI9Q
PNpHqvEQQg6MORnXrQ87K+MJHY7WZDyR06g6gJ8mJ+bhwqVlIodI34qwhMDLdQ3C
sBj0H3jBI1no6EYjzkISFmoXkXS4bOe94Si6ckmwW3wsOTdY30OqyXWjyXCy+Jku
by2STmM2nf1ZLsG/gVjoqzturkgQqwMEcis9Io6iRWSYbi1KADcPpjbIuhGjiJw+
6/kTR5SgJTir7X1vdM1UQFYi2tvIr3enscRAOjUp0r5F/i5pFr8+dGUQ4SV3F2XZ
i5h92nrJdsyG2cJc8Js6hyxRnI5Rkc/mlnzhn97U3SRrotifqtgwUE7+hNvDvTSx
8V0AnLyOoCW8Z6Xwy9yQbRC6WxMUPtw4TYcSaKmxabhD+3HIZ+yJR1JS3grdX11/
ahuXqiPMN+DRHsaeCJ7ye58BfUuH7JRvcC6h/Bq05gm9mYHN+ncXDpHMuB2mj3N9
H5fRBmi/6yx6DT8fDIJgddoCIKKCDXnkExp34PONUl3z0XoYZR42VDAiQ39ZNlnF
9VZ86DAAVY2GxghlyPLnq8j0pisrsRrNMHJ4jnULG2uEKM5suEHlwtKknyZZ/kpt
we5izvQfhMB7Vi2FK1i5N87meYD4t903UEq8UxI7E9McwlD65tLjNxEGxRMOFil/
yR+yC3GkxFl4NRUomC5UheiS5ikPK5FJWT7fykJ2WrYGRs0GursJ0HaEPnlCh2KF
zyoZigbM+h7f6O65NJs5f3wksceFRHc+4aXqGoo2N5cqHH6zv/Xk22zAnfSlMcGC
3TPBfVBxTjIaWu64hOmP/RNurqPiEQvYf8IleAJYzM6e6CVpSW2bSLL039/RDRcv
rzOM6MaSZvLDccpRL9LvkO5dmFJUOztrTZe4KizgH6weMSidgqL4E+X49vcEorFg
kt2QcV89Lqb98ehxlGnyakyTV9ne+xxVfonv358fuIxlpIFdxUsEnkqwDbbP2I5X
hLCGTzGPnrHs2sI5cAG1HfAQ3Rrm7DauBMrhekTd41EueuZdBLJypsmiSvrkCJk/
f9oF4WdP53ZlMv2HHl3TK2RJoSMF5pU0Ql8rwA3StsM1ltSsu3Ox3sTwjW69HC9b
hklvzPJJASTYZRHpinpCCUABaegNx9zKBl2m1DbI8uT5R55JPqHVfKnd3SupThYR
wOMhFKBC+4oYAU5MqyOQrFUa1QmQs8v1lG3ZBAOw0Y+XNPwWGCN8xi9QgSVlms54
EsWJT1FEsyD8vGHM9tioVNtSQ9w9BPNR28Ul+Zf1ib4hAEJ7AX23kd8T2meKrBzu
VU79UW2teFWMaVM/xkQC7UmFJuULiRLXl66RjEEJYOjxTP8Q2KffU2t9kP7OWKUc
uujnp6WliWUec76zcezrL298eXiYinhj9C00nzSDka3SBLlnnu/oJGx/CzrWAW/F
nctTfyZhYUKpnpv+iPL3SOEQPkqoZtMiir3b5VlgApgr4LDvdALOSBKXvYY094tB
TLLgdAHwbRFLBjRCB0D9Bbk7GEucrWOAcC2JCS5yORv2/7uNrqeybZQR8ZqT2sgv
t787i8h120hq4IaqGbtKPbnesvd+XtesBNeTeWYCTp3er1oGwHXnlpDtLSuMwcGf
FBWwqGdAyLfVJ1ouMVq7/YJ0+/FnYAyIkh1jvsiz6yfNMPwqS02ogpZ5yvY/VND1
SAWF95E1RNWZ5ywB7OAjq++zodIRWzvQ7qie4gFju7T6Yu4QCjDj2SHZVw2YLnEM
kxgNC+1RdKVFAaGajn2I5Gv9C2VCgeJ1cF2mxlW2FEZGQzLZqwTA6EyyP8l7VfSx
eXlgZr1A0SqpiGVNw91Pk4D9Q/ZAWAamkvb/PDRJ4FscqBm0MpRJtRe6u1LsTWLK
FR8eW5W+kUhoFr/cY+JQn9sA3hTwRBJwgftYZBeZfs6MfJ0CnecjTh7QNYsD6l7G
J7434KHKvDzGxSj/j72YTS61cJtbc5o6v+/URVY++7+RrOqbFh1ujHoZbiJoYGQh
SgKYTTWFb7V2RhV10ftAi2gU16qmLaiu44KpXfFuctw2Tm4pFGwfiX/jTbvXxVgG
DfpYckt8WdUzoH7Su1/7b260UsjxJmmNqw5lT3FXwEfUTu5UF9ASfn27yGmFWzXt
CFr4vk5k+YmL+Yr9hCvNSjp9Qae/WzTU9jX4x5epb6CY0Z/EjPVcx06BQbWE9JOc
yeqwFVCsyHqqOmxqZpYA6Z+ToYSIsHtaAOjCGqlkZxFSduGOSOkVw+fZSO/jTiy8
aRoSyorbt+utq4X/VYnk5rGeF7JLG1eIruaEXDuWwvtCZS273Z/DUcf0IJuEy21v
KBvyvpILmZTETh2Jfbfz2QRxSyWwY3bQiKsFykGk2mgrgiX3Dt7z+1uLtJqQlK2k
87x2rUSvcG27qkj3lGTSX/wkSI2/towtN1U6HHlza40q3RqMvbvZNTfdljzoYr/M
wNHIqUX+xFK6heIqjNCISUM4iTzBABwL0j/lPQOEo6u5yXUqZl5D3B11cpgbjdbh
NMpX/JBfQm0uRzbi/UNWvFgHk1iB/lhQe+5GvT02depKFIhA+LQ64nPfAAEYRhG6
eWPktEAY6k1xl+nf2BRB/6M8d9REx0EylmMzS/zrUOvGDViAcYsMcj2GAmbtNlYd
GlRI+K9l3/NA9MGDEjy5oE9caMfjt0g5XWNjtPsFH0Li+E+Uj8KxIXibtdW5Mxiz
8t2jHPrfj1o/tPBSJoMkB5zyRqlS5EBZhoEW4iUclmvuBpm0h2NuMPHGJeZKT62o
MFbkfgSKyCY3Cm4ec4c/ogQZkd4V/V4tBvfVoRyF52EBBXglp3seSsYFhx4lLsB/
C5CxY7B6t1aMpo2SzzSkh4FsC8BNoy+ptp64Rzu+9cyw+4Op+yznmXc3piTnF/b2
2gYJXnKnZi0IKJ3vrNjsr5r/QJn0MF8R8SKJf+jjZVMEdh6upCAos31AkjMXUZm+
rBRSO7pD/rNFKesJ27hZCI7whMAuaGg9Zwu0M5BdYKPbwA6jk5siVAcFnDw7tPd0
VvMbQcvUpgdNltprhY7Rmr8G17ZcH1mwV39cvELWRSGkIUYlnuB/2hlkXmf7IxLJ
C1xJCcHH4rbtupWEAJXZykprPlzrDAadk6ZNX1ChtFrN48PrqOidJb8U8xNF12Pj
G9aT7Aw+wEjoY6r4fx30tT+BECPbb5t5B//5Xno8gHQtAUarB5Ng0m1cDl3nHjVP
FvbTs2th+3eKxdCmmloxhduusJ92NDFrW1gBjShkSxVan5md8EFw5OTDifPZMt75
8G0qYGn8NalBjpsYhHx5jn6bWxzi/76Qo/dftHwEmS1avrst/P7SB44Y2/xXaZ/W
YZcMCXkSlU90jnYYNryqaC5md7/xUlCL+cScKzzvb0x/gCV14bYI6xNaPFkdljNy
PvHxHxzIqhDU6UAzdKEWQYBuqcvctpi/N1EWKzla6GQCSaY8X6FbkEi7aoxH51rY
l5G8jyDx9yJDwRp+SGMrFmD6dMQENP2THXFQe1h14LYMA8gqRIGqrtgNnSbd2YLV
8PFyDayvV7jzYYpt8LROMtrKVpdn2jvXfN3Y/SV6BBL4JQS5ZOcALZDG3/dMb1D4
c6eIwHki6plk5OEfEgZmnExzxeFCUHwsgu7/MDTrrAG3P6Lj+N75YLpA3Gu9JZGV
wYzd9RLvur0/QhVAtKm0Qj2DL7QlKYUNxJkM5sUBg5iqLHAeJK8uh1qhQYSxbbi5
olADd7KaLPX67VmsdpXyMQ3pd84nu54HP4ZVgDuRyCC2bqLvChe8sraviW7+z6l7
owhwqkuI5vNZXZu2HVyfW+xRVpYqtNnoj5ZpR2aoYf2e2djnlKte/JkM2+iBs7Xq
qtmHKhaDh3+3uSykm2tpS6LNjW0p0zOJe72pT6egOwEXcBpJ0GvyDwo3vSGbOFEW
5ukDEwJBbQqjzSM8GpySwaoV5hV4rtJEapLjoM2g1EvNgWbbeb+idbyMRc4os+TO
W09Rp+zQuvwLDGwmRReDgBlmM+3sVg+AtQADsAwEuThyBcOWdbEVqn1//wI+FAZA
4ibAhYy24RQCyapTducOECXFD28h8j6P+ErTJWXb45btNCsKPMkfuUA+i3859Yzf
kp+LPqBrUsPpJoEeYjLQ7ij4IbfPFJGcir49VAuZ6bcNxr9wrFG2m2Z59Ft2vy/o
jHMPsAyclXRrAMn+QjbiqLJFi07OAR6zKJuwKQGLjr5c2eSZM5Zpnf+Ue9lzAEnS
OasFlyQxGQH5g4EB/NvWQX1UfPsA8cBqRxKeDxyBsUnGpr6rWkJrkP58uQ2IBqzs
NJj2kUPcndAARevXRW8lqYMsG+hXjZjwwamRAA+MGJlRM0v7VJMIgAd18m/EBbjc
lS2DLw1Qpc717W+SQ85rLVOObrD3prRcgmT21MuBM8DRm0jZ40KNDfFdGe+CUe22
B46qKjx3Y4vdSMuPfqMimBYnHrFTqfoNES/ZRuu1OjzRhC2Swiv5W6WNfsw5zKf2
kB+6H6UB4MeM6nMQ0yRehXxttpVnmt3iGJPhbB1WOyaDt+QU9HZ/VIbiiClHbgU4
Oi2Qkj7FnFEqst3CvxrbiUfHUNEMqBZ/V1iYEv++lYemwaus5ZfgpjjQQGPENnoy
yLmUmwylP7vd9O4o/oB2OpTw2QwYLm+g330Tflc1zhM9fHWL3oBAg1zg0//yCTqa
aiVd67EAqj6BVgXNk5wN0lPxB4DaLAAMJTgJz0qvgsQDE37Na8fnJqEnlbDfnxJA
O3nDcWlfQObhhQJatFNilZc734nk/P+jJklYQPSJz80bVhwAtXfCcdUp7sgACi+h
+F3E8voGg8fadeMW9NnMIQqHUFHIAJxKL78jC9NMYLTEL8LFd2ONabVf9CP8IEcm
04Hpj6iHkU9FYtWgQwKtH/GvDjIMVswCjYp6QL31aG6Wj+h2iz8VbfsryhYBtvT+
X1vouFiyI0h9dtlZEIf6+lK/KU26+l+R5BhCAQG74RUQRELTWY+vG5QyAezdWxNF
pdQoPo8PmxpRUPGBPMqJPEDSuuIbkqRsGbGn8IIhazG6gXDWYN+uTiC903CeBUyL
JSpFBist1bzOgGWhyJTlpQ+PzFXWTspGUBaAYAq1aYnEqbt2jNgvD1SOZMI9SYN3
LepB0SWsPuxE0HzOehAPz9llZwAn85Flbj5MdfFfZHyQYhOfGptWi8GOQq9wAwrU
deXke8BHIN+ObQPtEhiP79wUqHAS9m4t785hKfJahO5NcXiPiBwX7TZaDb/w/JI9
cS0McDo5+bg6mxr4gHtEom7Xg8il2mUXUZ3AUHhc7YDPXOLuNGcdYGtqcT2TI3iV
trqIXXMVPgdXrVx/neNq13BVkRtwgVNHGzgkAv2nmLcFGienfjjalLUKrfiY9puH
/TL+awHxtxPHj2OBKDb3mZayFUj15Y4hciL0t6g2DpJP3nhU+wdx9prHBtQJO3Ln
TC3YXvtqB3hyVFOcsSFFdi82cRID5dfIjyiTVVeJ3yqv0hvhvfu+2ZTE8l9GnxLs
0F+vr9h7CgQe4VQ3MvsZnJ+PvgDwmAJFbjIDyUD6gBJHfyI4f8etY/Y7D/Q3cbmq
oCgMpRM9k0mRoUmNDVoOvPrcDa/csY45CeO+2UXJLalv9NPKpgF2arjPzU8HAhBs
hLDthzW0KOkzt9VU9kzUdAI8rZ9luZiTZcHPNHIaWmkLqQeTOLn4jgZt9NQ+UPDK
s6ak+O+4r8HYM5aR+FTS4DWdo2oi/0VZsoWrC7PefFwzd5Sod9sF915IizS2lsKb
YcL9qXk9ZzW4DnkALyKtASZXTDmz+L9KMXUIVhaDPHhpY8UhBXQPCRey24tcqce+
cSIK+uVYGUUReoDpA9NnpCxZ8pdT+Q2AKosC7ARel+Q093WuzxIzfbNeRxdzcisD
RWSzcRlQUSaSGJ/q6OrePqave7vNhn8J2dvCcAcJlRoz/5fQICSNiAyQ95Qjuqf1
A2+e2ACyBFvcMUCDlzbT9O+3kD4DppbT2Ka/J09cQVP3+B44PaI0M4hyz6F7QT73
XHQqGJ8ZTHP4VoNUt7Tr2cWj3SW8KpZVKSL7bUCGH14X2mESrNJI1Xk+hSZ8bj2G
5Aya9xXeGKVSDZ/XnDQ1kSdkDj2gZGHWn7mGxuttlGJKoP4lieO+XFV1iOH9Foht
OT/rex+h62FX/A1edwJ4fz1OARcanXvGaAF9BE11EdApXGR7rKZzeBqgPSj5fM52
/OccWtpauRSoYgbAcXAEnsHNpIBJ/YHV9jBxcZBCdYeXLn84XBfT2zSfL33QhW5w
8LPayQOKYTHNdM/fq4Lose5hdeiiXdg2PBa9mHPbvm7J2zlixzW4jNHRNuSULfYO
VPCQK0wtdH9d0zHRQd7FFjEwrcUPudGlCrIaQQxQBOc+f0ZyXShjE18aFKhpflv+
nxa0oTLJo+llSjR33h/FGEOAxsjAdLFDdN/ZVxcfvehN2qCd+wJz6cvcWkAQGeyS
zKf66q/1ifIgkNNuvHTczDJaYelwHJ49xWSevQmbaF/vXci4YIvbn2POVq+6i7Db
kCqxdQx/jupsTn2Z8Xfc8ztF8cbWqSbH3PEFgDtSiB5I90ZlpSlvKizPAGlx7uMI
/51nL6rbkdTr3BTcCYtxVU/oY7YL+uxsW5hQYl9uhtSH3OpR0ZjJTd13PBTwwr/L
CwiUVk6vQSfmFdQRx0PLzoN7zDL2FwBpe0S7m1Rp5UuwMLmmWdt+B0qYuQ/jWsX+
cSwWI0it8MnaAd6wYhHof1Azul5OmAZFXYBywUZekx71AcBQ1f/y0IYzf/sLTP48
Qt4o4L2a6jRXWG5ogrmE127LHdPtVg6jq4b3zE8wOJQlvfem99L3KvKxSHe+ccIT
2EazpMYCczZuztS1/i1oSaFesrXbmscXDKzlxx/Cp+4ioAKRwljv947a3RAlJ+bC
VNZ/4366k6fcqZXMIIt4V1pgNeV/uZcbhXHMDMBeB96vtUcFt+XU3gRaB7uwR0AA
YDdaDdAahex1tc7IAqJITHYfzSNCsFGPA/V2cAD6osmogDSXgEC3pRYLHJgBfD3z
CnzsjSjET/NAsQPbR71RSZQwwsLzMHI2V6tgXkfcIG2+RZcK7/gfm+ZJd/zc32qP
q+SnnnbKCO0CHXLRMw5GC1wGb5+xoMjp+wI784hPK/apOMzB7J9LML1nNbVcCZXW
gmt2y0GHXz+ODDANBytQdbiH8gY3LQ2WHAWMGvaUTXy5J1SGtWpufqZRet69OAm3
5NYpsokwyNyCkcyNuaHxHjMUbl2t7m8RyesVYmFTqCjFKZUa8eyobkWQ5tKO9lBq
o8HkqRVjg1y59ukbn51mhC91AV7qqf7EgKflory3dQk/QASdB/YgeTzq0JcFSMlq
9e6pVKVWTsM+DAIInzydFP/uOuh5A4dWmJlUdL4Die8VrS/2Wx7rDGNCjHP0D3sr
JUMw8BqpySEqkK2KukPm3SPs1rLjyG2IJYZi3hSaIRT9krW/EV2yc7or35WS60PP
ldt/5pOk4tmI8BXrvGUTbhwARCc793+H0QTYnVISu5YTFh+Gk+SweLFN0PJVYjuT
9bow+rLtPIsoEiddGjXSj5xcQQkZECZwbAdCgfeJA8IdAvv7DcdjOf79l/BKcizf
5VZF5o3bQwsi235loesnyuTix45TKKoVMHW5YOgnNhBc3VnNl1LgUu6kOdvQffh3
Y07jeoyd4OEP+MRotijHlqDLFj6f1a0IYI3C2sg+YBbIhYLR+gNx6YeeBTLZ5Y3l
4C2nGXVknh05sfnlWt33Hap5BUSWKyO6TM7CQ7RT/eCQ+xwmCZXMjLmYp8shMH+d
ttZtpVqbMUCNpM3ND1mqo/CR84gBMObd9N5MeG2a79ENpc9tKl1RE47RNe/7VzOh
UwQBusOmrHJDK6m0UfAj+NqAAzjpMnc9FJ+n90i8hJXoKahW+QNrMFDXgah1TFre
QSYypW/4xP2JuRw3O5puuULIfG3VlUka6ZmlLfW64CAi02SdDSwPkyf64H7B48aE
KwB3SszyLxrjEK/SfO86wElVvYE+tuN9tH4mqfROaodtdjvooVi/6drvIMQaamUJ
Kml7jGsYrhXzbOg51zAJd+gU8RaMckb1nExFX8OrLX5Ojk2OFfHZ8xqeVGn+0ERG
YsdHMm+5659kHBQH1vJ1zC+/4um3s6xC4BqMy9Ku2CXbeF6lf/4KUYeRR8W8MyaS
EJkSZ7KWnmYnTuvm0/StbfB9p/lMoJlUFFdd2BL5edBKGamqz5uI4PpPiYsGIzXe
gDRwWYOE+KnHNvI8xdPBT+ErHok1+BdHgr9w3moSfidhHYoNyM3exVR4amalV0j6
w+eoZxMHQt4zp7mXY/OUJHbxiZ6b5R8IjSTU9B++3yw53aui0oTDvrITlDarXlp2
uAkbdjt1JBVpWRxyDDV50L7MHkvYC53cd/IZf9qw4Rma7DaNKEng6vwjWaWqiOj/
MA55t9G9DmV0LvgNks83g6v3s2e1i3FkbHHXI7aEzgLb6rTf7IjE1MjGqfbP5P/f
/1oajW7WgIIA6kp0N+vxVCtN6PfiDB3TSpUtuQIUcpx7K51bVbhNdJ13yG3gOhRH
4po78RADnNgW81tWDFJTJqDAjYnIQ9jD+3vCefk6RAJVyK/DKxhcc71WGS29Hdhn
LvTk8J51dbOQ5N6yBbeGT1fwEliUBeHaDbULbeN9qmIF3i2FVk2K2H/HVA4LAI/a
aFjfB5WtGqubQbiTx9OlZmPDBieRQ38NAbnX6H65gZiHBCL2g12nBXdhc0yJ66BL
ChCeue5elGwNx2nCr5LZf5ZUgpxqKeynq55M663DLyJ+caaOLoDsc92pIZF0I1pe
nsa6f424mCg25laRywYhoZJt/o2yG2zEbL+fOm2sM/kHuDEECvYm/5aBWXwtP6D2
2FAE4uSvjKOLe2e+nQk/qfxyiFo6U/P0NOALDjJg+U3oPHgdBm18bejYPAzZbiO2
ToVceuawGiOhayoIIG/idEIPvwYGP3Rv21hDvQmh47uhYvEddjhtrauiVhHrCDum
v8hfuKSfFxVre+FKciI+6R88OIEagvUawwC8ZLwV5HXz0a10iHIEpCG9pX70gT0X
Nuq9LS7HYiXU+3/65HugWPaEvdCovbvuiQ33Z89NDm0lsi3fItoExrarqWHvbOKX
SPeQ+H2nvbAPNZg/uHnozjnZKg27CbcvX34xDRZVk4ehq+b+fRwEhclYUc4fpExy
AjqnCROAvlAfXJWeO1heJiCzaV6z23iKr29oYhGi3wZU0kCBHZC3vDwqfW6MvBqV
VtTA6s75vbdfAqYHmNcRS8VUUH0QWFoa5nnvGFz4f3d92dkgzccg/aot1A+rCAc9
PhuA2k5EgNvCNKZso6W04fa/MQsfLCrPaOgXzkYnioevzApEG8NmDenf8SVbXk2m
iifiqWI3rMPW+JthCzwzi8QjJdM5fuWo3BrwQx6MFoODs/aIFhbao6lpctG31LSP
S4m5yQCHT7qwh49ZWN1k3z1/oyT+cvF39Y1ejJq6inUdXbyg3ZPrZvor/T2P08dF
EStZFu0yDXghpbQIeCHLJIOM5cn/cWoV2MHFdpKUZxHxTSPpb67lMYPxAyaeMuBS
c1FJY5tK0KYNYXP2UkvRD1pWZEs0UpmHqV/CMaLi/bzfpTny+5blbtHS3685xqQr
Fqf5kpRWd3IZDxeBQrvyFPGB8IHECNGxI+mBLgGGazrxweqvz9vaVwgxYgEnYgxe
+FR76hjvrQM57hYMcLxNV88IT6lvt9Om1qtRR1DaM69Rr2/r68ChMMsnnp7Sw4zM
6BTNAdw7wcvJtH3WDscDWL4AoTeYXEm7LO7ITb0UDj4ER47fh0p6HnJLPv88V9/g
yrPcqrBpwoBirbVDRYf9ImvFApRuePG3Gera0aK/aIKmXB++L5DnNhL8Vv+hOobw
0RvHQT+ST1uL6zr4aR+iS79YFNYI+EuCPq4odRxDwwqGOdy7WETIyV22k0WqiqAt
12rG8/x3Cs+3f+Q3qQd93thqhtEPMkHq8/7B8XDrt5Lny1atXKn3oOtXP7sUCNWN
BjJ5z0OXAUwlrqH4gqWnbagloOOjnIwUG/f8nUcYL0C5QoRqhYpvcJYJuQkZzCzc
G1YV4f4yR+40vdJOzFJMc4GdmfyFXVyL7eTUUb9vUauedZaJCLA51XEkowLHhjYY
BtEUUCyqf8t+BRVYmkQEVo2Qiew1vFdVGdDDok9b0E4V3OqPgjzCzQBgG3xTUbwC
ml3dD7Nq9XlfzxX1IwqhqjeNrO/42yqTd+l4WZhg6Lqin8QssEY1O4zjzz0cjI4X
h9YjxATkFeKtYb8dlb80VyikWtP1vTlOYR18n94PGL5mHzul+tNv8QO7WqAWZiae
fld+dvvMUyXHs6yYoiwZiIve/Ab3b48A2siEsLGO9PCM5WYt87LYmaAZxxxezSkW
CTw5p2zdMWtuHfg67eRq2A7vRumR5vr0NjCw4PnWY3iaTPv5OeO9yAzx2g9i5eI7
YKARCUyYrgieJDm0adGweo2H7QsiATMQOcs3Ddy9LfWtKzZqSt3B42FZ5LyoVXwh
XGEBeQvxAi0hAVYIMqob+35L6fFYfV6GGlApKNliHjieT7ZEvZkcse4Fr1CScBem
4FxHP4APy3fK/9zrJGMCQaxW94Z19IE8DKWVC5l/nv2zqx8b7O+9eQXEUgQGnSjt
leeNCpXuswSDgJOPPGvz+vkolPkpwGrj8PT/upuxueusiHmjuhZ0RG23fs/Gpm/a
qD1AkmqXNz7QjSMFgi2q11beC4TT3i5T4gktHTR98WS90TfcrIBELP1tOg8PvUt9
Yu8BF/Ex9bV6aVQPa7S+ajdYUQsXyTT5H4ARYsotfka9eJlhelkPAm2e2+x/eFMq
craNQ7zweznKGDBsKeWr3Z6Ow1Luvl9Gk61qU/u/Ev+yfGD4vojGzeJWjP6yiH/N
fZ8wFNQSdWR785+Q5OFNZTHxIIm09VBFyBVn7cyqmusEGCHE3GT8NRIzvOYxuaSs
vqzKTGCj0i1xeNwaPnSG33MwqAkAiL/p04dWUQ55EKsVAhtqJVlQZtRIwaKaFElN
lqtLMIA+x3+CL995WxPPmWtKQyFTWVSYRodEcJkVrtXLNTchYLPDUAPOV/CLZcrq
cYUvLuxtzzwPlnRv10syUmqL/i7R9M94ljbB4cGyyv1oTrqK1fORwqs51YQ4PsHJ
u8wXE8YBIr1WYKxJJTr/SCHjwlXQ+hmUC44BEey2f0AYemHlBRP0la7HwWEmBgaN
DgVqyC5NsNuzZ2VVFDTzP+gn6GxnjSAnE+CL3ggTTYzZdUwwhOfzbnK41uww1lb3
yM8trBXmXM8RMp6/VZRjFxEJRNgnKcjFP2MKsLgmNdD88Td/NOv5VHCP/5jfCrMG
I6JH3spCNNWa9XHAJaA/L9y1KdjOkMCqliw1ChpcAbkyMiSUYqTthM7JOIicwpJx
J3PWqaiPX0Z9AqKEvxiiccd+LHXiet2jbAn00IoK83litHjDVkwAT96CWyvpqIH+
vREZGhKICz9vzID/2QHjQ8qlEv9AuYN9FDNwMfv+RRhabFP/4b2vj5O+k/OmYphJ
lsGof+9SxK9wonSeY96QuWGLC5ItbfnAFEFiZoxMA6chOcNQk21Fq5RagjRQyTM7
qjyj/BBg6mtuOJfWP71EhGf7/QaeD6ExcjDsO8ytWgImf+SGHEQMyMwkmZcGp8Fj
V7u+B5BGurfF1g5RUfMYa59t6VM3iHqYBbm56aa7FSmsAXSzTUa5g3HgF4ccVlFg
/dGmcX61JfNUW6uqfrZ2XZtv6tx04zmHcqR6DneuGWh4PyYxnR3RUyCl/c0T2Y1T
SucTTPQU6r3rIhxY2tQovYbfHQW5fB9V0aCNArYXVfvRWY93ERJXVJe+4mM/iz4v
x4BXR8k2gSudiEuvMdOQm3sdpqHUZoyTUWAm8wGRZhKUN3u77W2SSx5ZDgUVArQ0
lTqM5cgmIxcjFAyH1uVJV+p9+b/BnR++uEpw6VRdiGaCR8T3XjiJNhdQMwWnUu3q
LZLoLefWk12/6bcN/madwgab+aaJsmfDwJRoqbfxhz3iYFpaDtuRaeK5NwGR2t+c
QaDs+NGI7W4F2rp0wwABJB4lmFWAmophOc3cfbtT19ZZbFayGXDK21eNFHZ+T5bs
11nFwYIRqzULFeOIIz6ZFLpHJq2yTPc8aoEgumqCdKDVFXfnJjhCUPd8wFCCyuAe
O/fv/9msBHpc7ULYKsHxXFJCx6hmG94qaAF0LEkQrFV8iPA/iCtD6+bCCkrl0sFw
aZIY79/0EMEkV9Cvfg7bNWJz6NFueq7HYJA+L3iQxrflgGk5H4G4+03UJLWZa5ht
9/RZBnvM3r3SJO+2Cv4rQjKxWeuZpzt2rrlBlpGLigobgEcqN55i+/gWS142ulq4
jsKjKF8ML5mcFgPawxyTXx6xHvwklhoIBHFLYORMlDGgM8ObHo6v+bm85EnPSkax
91eQQT3URvxP4sDwwGM0IkvFG84oEBfZEcX1nNPaAD9MX+s+9J1huwftJAFXXaq2
vc4cowWfHOKCZv/SRXLuHeHJKwKFW/0V4F1Z5ltHCbJO5lvIsfd763yvHpqq8EAy
gB8GVfpLZ6LatkkcPvV6/GeUxQJMDxC8B9NV650nLiQbOFRKRzzbcaZ4RhSe3lbL
bgbSUnysm/ITtms9/HNSQgWiIzSsFo1FhIHmzeX6SucjVZXQRZC0YqOM1hltKFuO
Jt/yYAL3GGJs9M2yFkZ5LFOC8m0jokUEEl3ZyWlq2mjqGXQEzqB2LHrKjNEio2jB
qZ1LIZkj/UQnNH2caLZGY167RzSsyHAtkgyVwSLDkZoziBKpMP3sx3X/6GlRpd6w
7u5MAIiI84IneOOK3cFgQMfMJaiKFt/RuZY7F659jIYgwCgNp/JUkXdByBlx14fA
bFEeJmlSDSH7Zj6llk7nGHnSwWdTGUnqURNbi9YPE720F/SAH9UhA7HfdWQOEA6c
ey+U/1XqZxwJ5eivE5w9AIUwlUvXV1szGujjryX0fJuP+BOi6upWxKc78hFvaO4j
h3K0B0s4GaO1siKBbb+ffiHvJek+KePGl5mVNnofUHls8ofTwGEPnPnSWPeN4K0k
72L4oMdKHAdufQLMbveK7YRjRtb1SFXrym9UZhUo2aglG3VG6VecXKjxbsdabszq
HNV0OXvKggU3nj6Jf7ZPiD5HNuS993vmzmIJTq3YwjWLbf6ecNAF0tRBp2KSbTDa
HXrRNWfouldsbd+++OtNiU7DNuoqmogDIEEiiCbQ57YTcNtzkjkIsatjwfa3SGrn
pf2Sd60o8k5XeATthJQtywj5ZJNdlXNKXFczuwJ1eR6wldzmc480c03gjnOIku2C
8qQBLtzSWyt7cwdbmwF24i/f6x6LI5Qwb2kFpS/EqSDBuiLmStJEciFcp2SLZ4EK
1JboX6aZzByXoqzFxHwk97nPLlCQyaGzF904y7uvvOya3IUwt9uHMUu5E4ZPfFq2
JS7RPqvDhv5joXrfBX0eAFzg0660K+P4F3T7qIsE4DcS2rY7xEA81kN9T93q4+Up
6kMwswWJxZU8mmZjGZ8RTilJ4DaeFDZfXo4auZ+WlClNMqH7eZvdEPSSndY7Iq7k
NsH0R8NmQFHHhyAiqXnMQz6FShxGho7SK1/6hKCDA4PWhjooPhOp5BWMcI+VrH9l
0W+N1CJMgZ4drJkIQJxZznQ6U5i6QIbHrYl34XEDKunNX9e7FpjmmgUIftZgrMEk
5x0wMLssnf+lp0fOHcGsVjDHoxXmkqySXcohc/7fyeNrevaZaWRLm59e2xnecdVb
/KmcWtJ5vYk67hNsyyWRDzQFhNrZKLkvgMz2xKoDnWNQgZU4o8xN9Ofb2/AVgRG9
yVyPx/ZSfuG6xcd1ZfHlTn6zcBwRQAdTI5lOXTnHCmWuhzAyMHW4F+UFONCuDVm5
KhnJRp88TLNC6cz7+nJ2yi4dxfdTqHscxoc+aZ7bI3yZoH+FOAvI2M9w4SbmEZ+c
Iq9jHLUMI5UVwpV88EoC4Du02LvOE+5st9H9TrfoDQiGJAg9906VK41Q/fH0xJvr
u6uZvcep0iXXK6iMlrcz2L9Y7LIQzGBtWhRH7zC4qnfCnNYSae9HLVS6e+AJLxiV
uNdpcDPwo6cSdciC6A6P7Y9LjQFJxgpymR5/d5JMiSzXHCDlflKyVc/Lod6TClqA
1kZ26HwQQlA4IpuGJaeq4m3Hou9gqQF/i1Fohn3XwB6bD+Az0LZfqRNgoA4hx/H9
kanjc6I9VHAveD5XZvVsEKxmSKj0CZqm3h+f6KQlkpJS0o0JNDYmHmt3eyOFFfGu
iFUlRwtNcHWUmGH4yG06qx/PpNYuIntd8xz4BTQdMYGlc8KAtc6Ex5xLN+ztCU4w
515uvaKkPkwuQX4YO3DrAHQcTousW3wdHUjZ/1Xn0645hOKwfwc39tC2r7yHs6ro
1Lfw6FxUmdW+4fmxrp71374nWYqqkju4gUdB4r6/E9iWCjHVu71z5YHo0QU20r5S
2UL7+IETY24zul4Gz7Aha4ztDPD2fuz/mtSAiOvBujrxet8yKY1SkUtRJgtK/5V6
CpMALqpWr8AqG/yUXnaXvcXadvBRlNrdbPhnPLenWLEIRGxz83pLaUEOi7i1O8aL
h8tFUuLJ+9BYP7JrbkmRTr/iBSxcZ0K4oq01qyiZFMcyN8vvwlvvtauB38X4yHiv
o/XX7cQrgQVmqbovSi6fv/usBRAJdBT6vUX8JSK6+2IYqD4BdqyyLfQb8PUWMT6R
e31+pzpECI4vFTG56ILV9ADpnSakiBEDLGaxGERM8co9yE1szhAj0e3EQiDnmEg2
thlTzFpMPdWLZ5mQObNU720yPhvyyJOLlsQI+3KvSUim/Rw8vZfKZ9f3VAZZaIAV
Ou3jyRZuCoRWkjyNNAAU6Uo03kEsZpltakT7jL9iQ0/7BERjhpQUFNmzoNb0gu9Y
CSsFlmuFnO7ysNMkZUtAsgZ62ZtSFQ3aLs+wJQAYq4a9+rgL8QUjyHWKay0ba9os
I4XIuITbnruyiV+v0fFKCb/FjqyZf25dDLCa3YeVoqoVzXfIoULB6f4nsTcpE/As
5I/s/Cnp5eEzThqVFOiA9MqdMZaYZf8bmANUEJb6OVB4uqMrrFkWjooBTQ/r9TXu
SkThgLhy+zn42LpkO3oE1mOmK3CfiWhYgUc6+xdAOzT7sMR3x8yiARAmySyY7OOl
SuWtwsWZFrdyFiFkXC518P2J18MSU/p6CTbnS5XImOew0GQPuZlhAvZdG7heqeGF
FvfpkhwH9ZDPjha8RZ66Z174KGQSX8VMVhVjSZdSqkce9gyNaEjzwN2kFmzB3voL
TiVasmAh4iKOXXMpMqwKWVygn+jqJqtea1JsXu6z2jGAepVpqnaxUldh2KpnqKkG
+yWY1yUAd7Vt3eip8QNJADF7jFTff5dXNIvJymlT+X87+LjSfMEvTPu4PSlEL8Rz
HX7/NXpK/sm4m3301o+K/V6ZToAP83xq3qVWkTGoScA/lUJp2A+PpNn8rprSBVyA
/po0f7bcnVLi1shfb3nNnrV/I7/uG2pIR1YfMvzOVfbqmrX5K4IFT+5Ia3+X3BdV
pi3Yb5JsaBV+ZEImSCgl7nBQDOnGV41bsao73mMFlEB0taVoH2qUouvUq+GZ6lco
9l8j7wvv5CKlzQNvV73UwMMvqRAxitAyOu73BUa7NDXv6z1yxWYIGco9+MVE/FiB
Qv0GwJLv4VQhO8g/dQrgeKCRvNrFtCtaQ3qACH2XRUbHAKXIDgfED50xz4Jd+Zzp
7egaWa9MU96WlrsJcSwkydBTb7fDbmUz5cDG4lCgg3Z7s6q4W/3vHvvXMD0pdRZn
0wxV9XawIBMlQggPMeuTFK3nU+YQ9vTpKH0FCtjnB8XroZEIgoO1w3BlVRT/1dY/
GWp3aaQoj2zv2Riu0OcV7jo/2KAVf5I2ME89mG2jP694C2AUMs24OgWVTxHY0hZD
ooAuKHdRXuUZfklOnTDq+JL+9y3YujQZxEaJ9ahXcBUsAT3FuRkffxVEO/1Mp+LR
+qHCPD//Q11dOfbITQyB0e/cRNOvgbFrwTuCI1ASYGWfNoAw33OmRyQVFcvznTMU
N4NJ+OkxRb4NQ71lm0IxDkgufCLpiCKjdEEzSAN1Y1lz9YbGGofn52kad3gyWuG9
wH/baDoSYVsPJm570eq+wR2kVeADaqUfDoZy+9E7Drz7zPFubfp1uJcaSe75lSKg
jy+kLNGOj6jk0+b97w959qDO0RPx3QiK8glOQ7fIogFMsobDhJMluDheMDrTgI2S
Bm2KWN00Ato9inIoH9Xs5yDz6N85qhVl9mLnHHo18meQgV6Blnhb2UHVZ0J5jgu1
iS/1FQNLWiqOXs8+bkL9zzBGU6cQeuTtrrbOtMauyoomybT3ANzm/EzeoX38PFQf
pZCnSPMPLJabSmREFkmSX1TraTGgD5i/myapGyikuwDfmZCYSMiikqVoroIOCorz
zrcevta4xNKIF7zAG221C4SOPJYLvu5akooQiFo94ZvtDFdMbWceezbsFNPq2UE7
nH9NwrqzrS+SaMPAOAq7amLyklWeAHz+JmUnrnjfM2r/gTU/7+A/Ka9wU2SFTEBn
DR0chv5I4QT/a7dBCeI7njzEJ+2j58+1laDrDviK73gQk3N2970CZ4gPJfvDYxCt
zViDwsDCUNoMYcuxqehq8tiWjbT+xlcXIW3xfnntRfXCEakPFDQxub42lrs9mn+K
ftQMXXNhuQxDxAZLOfJKT/QyKBsiVvcPbyGe+A8dwCUfOa5B5/mlSqxSItEajPiL
+ufS7n72VLmmxRVeM7eY1DPqJw5aqFKbPvgQXpiJ8zv6mgzQW5VqjFru0X0ze+Z4
Ww05dFx7hpRd2nsjOo6ER0fMXt6QGGqc8ji3CpI/NoU0VCQ9WF3r3Sgndbum8mMq
mMF7xUxce48fPhA26I3OJYBB0MeKCMpG/+Q8SUxc93YkkRbIocnAVm2JLIDMU+bI
B+CP/AXZXktjUi/Lz6l4sERwo8uL/7fdulFTKVwJ859Ih6Sfecpx7F2haWtWEqEQ
DFeZWMoklAjRJoeqkLVCsmKQySqx6XmAC1HCqPbPc7oaPkrAUMDtHdJs1XOPobaX
8/FoXkQK1Imam9/63nk6ElFQSsvJQV9rt8U7cowmEBT+VkKj63x+i/7o6JJvwEkR
h7tykmBLsmcwWQSd0EXcfsv8CYS5H9solf+XLwMvaCGN4ff8MrBffio/s2oUV65H
QJ8mNI7+ubDYABvix/IicHYBTerRLjOWMsxWcqOHaw3B55F81AHTUONwKxuVDOuU
MNazG0qrQn7gt5SKrQgTOTWzyAHN/4M/Dz4GV0LvOyHJHFD74DfcJVnHtazYik6I
su/M/N91HNiD9ud0UK90Ik/YClKmrGBT8f861CTmTlfYHbAdTKCCjEgKOce4ZU8F
/jdY6O/ulkr79ig4aW8LYp41uq000WKiYn0tuDn/AKj4kZmRydGDBc0eZttMCC4E
l1p711p7GgqEY1SfptLrHXUU+cRDSPCLy9ilwLvukEYiJz04nADwFohhZj3/X02Y
+8VSMgoqd3lsA1yyvXC9d9/Xnqrk7zkxzw8n1ny6B1HnYObm5gRqcHSSd7B2srS1
nyhxXKLLC1nU5BLrP+QYbvj/62YbqV8WgKmkXV95Kp4Xbza+ynz7d1C7kor+szC2
0S5bfBKNLalIVjQeDlCFz7n/qwVkIzSpT30ILchzPeyR3pZgO8eAeIxyoDODY8wI
p3tpeliNobFoFj4jY2IT0dQ0mWgnpmVMbj9kJXLeK/PO2b6WrVXb56SJR2U1aVmj
RhnH2XsXIJjJ4ke9qA+/BSd3T2LN7pLTA54NBEUsdwmEjKI/ZfNONKNQm90Hoz5r
mvizR9eu8B4WWFLerdIEVcpB+mefo/Y4nQwvoAjokQwEL7VXVpC2Acs/vxRwX2fM
g1niqlotTvMEGs88oZAgNlXbUuAnhPZyrqqRTKm1ehiyeyda1BYlKbihBNlo7uAj
ItKGD+7RxeTA0ZksPouLOnupv4rN5KipWXU9isz/4cW8P1ys6lYgqPQUfbYEbscF
9iaQqC+L0m3gJ4giqwG73OCwOMHcrmcOdRGd5FNgzO04gfGZ7y+IDOR4rs3al7x4
lGrn24myC9PnlZmtJENkC0b9yYV/f6BaeL4eQsf7lWNykvW6cdtDnL/nqJHJUmKj
+4WpWMrp8Z/3IrX4QInEk2L+y3WPp4mbTpNmFEBG0tHviPssKUDJMWIczR42kcHd
EwjFtn2iQbAoXKCRmmJgbShfYTKZwNbjphf/sKW7WMLPwP9i3pGaxwcbsdtkk2/g
vRpSeB3P+F4d/SvHtYZCzVw46lV309Z+2daHzWXxgM9OY594fMYh43bv8m3bHLBK
L85flw3vNHHW+iLDti2TaZDWWCJeVdn2e/y+Xxtb0+/4VZ0fK6a4DkoqATld56Vr
0KK3NUt3ASQFHTbgC+CMWnqqGKbzv0VshyVJy21sgnSdFFuaMCNXCu+eB9ZcQdK3
GoKkgMWpTz0aFt3MjuqdDS9TzqQ8SMQsbJK07KLiZiUW/EAnyR7XvvpGcwwuRlfO
r94eLj0pMeobs26sK0Gjh0f/US0G90lUR4qWqMufV1QffvPmyg5WYc3Bi4PFEJHG
pRKIrmdYK0goWUIH0Tt3WkvZw6HX5sETliN8aXE5TqYa5ZBJWtUEIr5HBdFZoZ4O
As7tthWXh1y/ijj5udWRFght8Ji730uYH5T/hWJ16Of9v73MP1Z1v7a6kwUCEKgy
CyMaZzDJikEbrKBKWHdc6d7J5Ntt8DKyhHTVaQOyN9OttbwBQLwuV0OcVgjXw+dq
ZOfiLvDFnx5uC/c3mAjwjesKthDeJEFQexOqyfYpSJeZLpuvrCnh54SDbQcJdTjG
37zM6Mlg611NJ82x0RXH7JAA/PFx7rqAyeRHlfRklgu0jy6ejTJJweQTKS/t8DFa
JpyXLRhaJe3rGo5OxXwPyswRFdjzsfUuZFZ/qVQRjdNUtoM4LBOir7aAtC6QRsuI
EJeQZaG5bn1b7FUhjWsv+EUa69CK7/D1Yri8MQBqphs9fXuMQaK8Vt4/wI6miINr
J76wNgMU+GnKQcQJ0v38LR8afcQ2hjbtIojhbKgXAkFkkEi3QTi6shx4kRjPehvp
4jVYQ4roP507jDDAtQ+OQSh7EQj1W9BojXEDNPCxsEWoF6jZ0aU6uKTU6TCsrGxX
Ul5wEhhn42bb2jUHdlo+SxYa2tqnBwPBj4E9QWwY+6nSWFbTmCD0R4dJtbizksak
zBRrx9xmly6eWHF07k7WxBG7xef6YJU1fEh6S/mPftUmQCX/pnSXpoEZOEUdIatf
99vEQuWHozheQ4xTMJe7IwveWvEJ7LlavXROKZHfTSk8jWQULiuU8LgtYw6ZhXFg
pNcSs4eKXGIODKLkxPdwRM6ptua+EjQMS9xZqo6UI0lGqU+T6uaAwVVB6b30CYsq
Rqk/XOPxUbqDjBkGaWTNvWcRj0roLfGZJFfcwLWElo/hs9RT22sfprcOehMn4KrE
C/aIoSkJ/pqlWDsp82dJH3gVIgC9MbkqRXfsfmVm6MWQDFx/SSitEFJnItuL5mqM
lzJvrqFHFMFS6XuAGyn/EjRWki75lLC7VTjuMHZEn1h6bxQxBtxyUvuW0WqCKNMc
64Y4DKJbHXF9QscbvWOzRaCvUo/HH3JJOb4V/l7gLXq0JuV6ci/eZVTly3caKMfl
c+V4O3Fj5jJGOcf7HDiZ24GzFzwz/ZS6xHvyPa7A40cbG4FHtVAcN3NKpfOaPPkn
Duc6gPV4beERirGj7iMUXheArwkuzSsxsLLINxq1wVcLWi+7hGBP5yE5PWrBfhA0
/gGWS8FJqqs/ONNZgBCMNCecRBZwZJ2oXVC6I5YsIISFzgBYs+TEJUVL1Q78xiLO
wZB4F2NWawawVSauVVawCCr2JCCVQp+zOB0C75DlNtEQs3dptLXm/FsFhH9eyvJB
3ElbmuUPUTekdahkHPiLlWNyYjVkqBkjYoG7CXPaRbS8zBWKT7Ut0tAWc0oIZPm7
NZZnX+as6B826/3eeIkkpHeB3/bcbP4k9CeFwctlx9rtZztaQHvioW4ae1kBcVxy
W64aENPXH2xe7tqZL5ypHBzY4ay/KW++Ybyk03b+tWJ+TLZ+j3nyeKoN2FNKa+X0
cqGK0EIMN/RIjIsQbKPjbnmCqAPkY6X+4fMPxd4FBSK2umI2GLzJ8uwn4+rT/t9T
64OhhdNDsVJZrpmtkwOdldXlaAkzXP6nimZekoP4Q2IKpbAGmhSImyyJiRqZUzQ1
pzkFHAG/sGlSGTyBViL8d4CipML6fPpBm3RSZx8Aug9VCsrAXMAkuYXY5V9m47hn
me4MJPc7kHURvmdVzEi+3U86S8c/RIZzErYgkpN1mm4ORAOFb2yxnumbbqca98F9
KIitCMw9OCvFYBAYxaeAvQCyB9/8NWnI23iPCwZmFdFbv0Mjmr2peLS+g2RAUJfb
TPBne4lu/jNgiSxnsWUCaaQlu4wN+qBtYsyDsgLEAQNiVx2dJYxHoaJ3XfVbWbi/
NiZKZDoqyqM3NSzcvskkBYNGNqN94KorNwCkt6eG74CQsYh8hX/WKsIDkgjzrnDk
LOOFm0I4bqiMcTitlpMGILJRua7XuXmUe8QjMqDDX9ELhabdh+Ry4zDu4FcgXLwm
dy0HZL28IiXzHVxMzAXopTWVIFfb8Ub7+vTebJJa19tHzt5WrIa5NdrDTXvMU84Q
4RVHS59IDjr6CiZua0UAUHcQSmY9Sj454+pUdOnPOgXpkgkkQx2mHy6SfuNc9h4Q
Pwemjym2hjR+qVtH6/YOm7F7tJduw+Gb1yY1Ab/pYgKbP6lk1jq6g9mVfpUYPZrH
x+b0Lc4QJHKflz82jGx35F4unKQaOF60VZ09q8DcQGVmya4AyrhEl9GvsrxnyIdf
tpGFIxyNLgYWqh/9XWCAy9tpP153LPtvVZu/qpElT6rTMtSOedrTCqEcc9XYJKaH
KCfnoPox45eBnrAmCnYy15DROuncns8Ba4duztHabcUSTT9a4ViQ/ZLxlVQJ1iCc
LZeN+et7EyVrXyDC3afzSSp6KCAIKksLuXooEdByexeQPWLM3IZVeS+V+gV6Cs3N
n3DYQh9DnAZbIwT8BMpfX2SB8sqzFWpd7KTraVbN1W/rZfyDka+++YC7n8FZlELI
jym1sUADcawrt3BqoKe7flNxDpUr+vDbNa22hJzd3WGpXRvV/C6RILqmR1nmSn4k
Q4Grg3RKR+wbbRERDvfqqYN2qviN7vTs0uH9Cb5v8tq9cWpFL/bkN9ScfC0dw16g
7r4ccbiHmTixwEhsausLKvIYv5EUE1PYd3Ts1ju1ADMtp55YKXKSG/I57FZB8gOl
ZtG+lSHQnyvpsN6YZFsQBxQ8UshbrbkZN4W8eWRUPoCZTLTBgHHdWN7hWXJVAvH3
3VmWUQg2QQTxLIIREN0Mnx+Du87QqeWuGiqV0KziQigUXnwlTGlM9lQKLd6fwkJL
QQxSH3omKbAy3aTEKkwCo1jhfyAuzy1YuR+YsEhfO4CrnoiVBebtgB85os2fM7H0
M/0Yz/b8nKSDk/v8T0v5yKhOrFYf9kLV2ycvkioqMZeYvwvFiR1P9a5NdxBmCo57
HsVUmnYbxNrIrl35jCmVAiGp5yqsCp+nv0kLNgNnvKOxGopx/GbrCutEHEbK/NLk
XlMaQM8AGIsEck4Wdex7kuvkeFChQq57Tyc1yUP4al2vGaLiV6CwoqQHFE4Xc7a+
5C6JnFeW4iZyCUen2LSryBOAaphtsGuroxoPKCUjRG+k3CzrwNnpYCmXQJcj+sbB
bxYnCYnWVGpr1h1YoyXPqqax8M6NAjH2Fy6XvvfDWESMs6AAvvbjzeXptxSaq5wm
d2q1f0A3SUoqqcbmdq9c/oSKCu9/DmYNW68Ym7+DNHmRFGpbM/EQ23lqZRIUNd0B
hYZwMloYp9vp3QKPZSyzms9lBQfmxHLvAJ3v/JamwA2gzfYdBJL79fsWrqlPNAqd
6iCQ8W3olaUVO3A9/IeQbLbXn7pK5VLR3lmxvAsbmIBZOMX3DptZYQR1p65RrHvD
hnAeZJLYRIwG5OIcP/xTnDkhGt271wv5CTFaJ5GMeL79p9bJmJnOMjjMuk8rqPAE
7CYthtQjcDqdGp/QzkrILTKN5igxDmwcxKdAjp7JzxLfUtQplOD8gp68fC/9fcqj
JdPYd4O08g6YrpJgfCuRA+rvCAjGJZ7xiNoxV5Jos/V5fN+OxUhhXFvwKssTjh8W
gZq80B2UIzfhhhWcYwWYpdVyEZ+EUOXIsCMAOufeKYoJY8JDB62VnB5zG4BQWw3C
J4vTq5btCOrsvVT6ONlQVc7IatKtUKQW0j7H/PgghkBo9X8A4Og72h9r0bj4LLCW
13WG9wojsUy9WXPzEIoqWAGb9SXv//eQf4vVQubmDTm8rsymp4fth5HoFMGp8sU7
ih0Pe0pKomz4nzNlO1eAQs4OUagSauYg2PbLBOnDQbacAf30dL+7tV0F2fLmAvlb
E0zFtoTEQe+VVMWPnWRoqpYj3qeiWWW/2ANt+njvxUS5fcofc5Cx9Rj9g1K66IRd
kLBxzghZHQ8qr/+uvfl5B8fdXDmayXCC3dkWYPGCNWjCXAjDxgVhWLIKi0AZdVDr
KWQebk9SRQ2ka4OvWmqCAW9lvLEScXGa4GvXNLrGeFFnGo4vx855d7YV4Nmh0oeR
jv7v1kZ5EVeZQeho1dWHSKOfUaDU5En1fqBy8nj+uzsr1KbQnbaV+nlQa8OPd7t/
vjvPwsmuv4fvplvFjipxzHhQFZZMnF99Gc1JaCqvy0CTyVSqSOPdB2M5vj7DGLJ8
unT0ZEcrVcbFJyu87HkGawZ3a5qRz++M5jui3kjtDldiDZnO27fr8RZFmkNBWAnl
elmtAYjfI0myOA/klBz+/4bWVe4IaE7i1ksT00T1UilYBgu6qkzCE6LulCzjNls4
S3T5ktH1dgAhjUs6nJiQ15G6sjoY27pN3dx6dAIdLJ8JonJdylYF/uLESy8Jj5jg
34eI4yf3xjofIrNmZbKH23/50/onQJhFUFmmc/r4HVyvamWNOBRxde/XU/IwXN+J
s8/HN6SaRpqyD8ZBjUISnt/Lh+yEST8kEiSENrmnw4Q1B/MwmayZpJLiQ4bNvx/F
Q1MK8vE6DIVWBtYjGdu6jZt/OceWRFIze98bePlMPdEAZ33E4YFCFDCW/kF4Z84/
lRcCpXOXg4KZ49/6YA40Qsul/j6x9RdzX1B305OnWbgWObhvc1LNJwVdEAvslVq4
AVvLBkNgtibEzD0x+28HHzYspOZxy8r3iF5ZjWcScMWfJgpSU5V5P7xm9sJr35aN
yGvFEJHrvUE7U0Kme0eHOtluuxq8G7VAIaSZH8o51C66ODrLx6AjlOMImUT6Vx5U
KDmZLSCA6UzyAbk/laEJi0XO8dBcoMrVIRrlGgF54mzGblaFuaC2/rtj7wdHiey7
zQQYO8Q1IkAqKub7Znga/CtJVQ0O7J6Xoy1hy1tlU4wPkC4caHULiBl+Ik2nO7uK
50jjPoC+LY1Rw+7ycTwouF5SfbXJxXl9oVOmHjMoiUgFDRzHlz158mhRGfkXd/ki
3LBGdgErW2Ra9CGqzBonsFKGHHAa0NOnjQvgijXzNuYH2reqbSaDKC12bbVCTC2L
Glkhi7s9ghVO3fsNh58hB6pIXFtkuXGqDNjcAq89pk5uJ6U3meAInmlx+t1QQ5tv
oFvvzTPcMLf6+BOmT10q0eHmSSXZ5SH1IUrswxk7VBRVBPpvOLFgab5n6ajDyFIV
QSgZLI4WsM8xsoqHk8tjc28pAxv2oNO4/zeRozJvy3TlECuAuQm23TGam04Hcsok
1xrN/fcmnWRiXEyUecKLYA88xBXEA+Ief1yRYdsMEnDjXF5PLj/Dk839axE5Rhlq
E8p0Yionz235RNmk9x+mQwlAMvXIQYmg8PRKtoEytcWHzRwdyYa0lcWr5t2IPXJe
mcRIhk3RiMIMNSjeH3S5WK4oudZi12yFUE+eQ1jAuWuuJMskvQD9gicUH2NC7BAZ
2x0xMIaE9XQmAy9Z+Ob+0305p9vjBVHG3H4m19Jkv9KnFIVVUFljM7ktPEXlfk5Z
Fvs1NN8CyrMlH2XVX2H+E4iX79nhQFcUFOQ09yiiy5Rda9o5nyP3uFEwzwcz3p+1
6wipFfo0k6ByD2ig1jkc+SFGylYO7IA8SYflXc7r9Oy9SsL9UAxEJqeQ9SSYN6yU
iM+MxRJHrNQRkqvjnL6gemxlMKc4fxlB2GhktQRixT1TI7cMYtpEdB/wvcPR/mp/
wHsYnvjPeTr0S70WdZTlrEPOcXGdgeA7TfNEXJcDj3cCLaewNlbfUGPkllFZjBeM
1Lg3StP8ic6s8Ga+IT9SKgPpNEwM0bsTZ2NaEzrM1ilKjJ5WnjySWtlxyMROp8Te
cqWPQhEmatczWlNHUFoo/k5jq/8BRmA39A/BPx+sGmQt0egldSop3uYtKQPTE14p
B33ytC2sRHJpcA5RGbHA+i8rR2Pd5Em3OqUn/WR+mp0B9OpmblbK8WzkHxxuZDJK
8XG/fAsZ+T2+O4U64oJJ7GAvyTsj6z5w85O2aVLUq0Jk8x7y/OhebrpkRNVnQZsf
SyHFg5Bvl94zTNl5qvwUVmEsf47qIL/YT27q9xUJOt2lSV+1h2SRbCcBa9dS92pf
71aoGAmqWzUy3lGiPPnayrHXul4T9O4mU/4MSaUQsh79xUKwLgK72OxHwt4Svb1U
hrpzvReZ7WWrDnu9fyzt2Xg4LeN2/S9r2rqAwaNfTL4+8y2XSLJU7YXFQzB+S39E
XBMWncpIogjqVipRbBYIjUsBg/lvriqkUJUrCCYXeLbyUAdrqKBgeDe6vyygSqyp
+EEzv80ExXV3nIT4Rvx4gX8q/jMkLxvtluC03i/FDLrTYdMOyOR7HS8NwN4CQfjU
Eiq5Hs/OmUvOadrte00tRiWI5QDwS7K7ut62Zfazc+ykIcHC0GG1MzzzFMyui23c
v9Ttj+IUAC3cy/LrhzppedbMKIacUmBTdJWxAoizqc0FjVq2E7g8+8tQQJXe0wnH
MRDGci6BCRUNqp2ONUUBUozq8pjFOYQH88XKXr/m31O92z+TWNAh1mE7zbb0WvkL
wQ/KWDloAfWip41kh7/qToszQKq26m7J/IXAJntkVbaahi3RyMXq8me3C35rL/qi
zq4z+IJ3iMowlfBEVvPZTWwvu+s9Ewx+rGQ4J8fu/zCccYMruqXHej2ikTGw/8uz
HaXCTskdUI1uFy5pVE8VD1qsKDPtUhreo7gmUQdAsM/s6Yttw/Om4RAZJbseG7le
foIRIaCwxinwro2kPxnL6dRFbP0EpNOOTW04S8f0VL6J0iMsyNCl11Db6NKnt0Qg
2grb4WzxxTXw9abs1usAJ1tEtwpkEb/Xvhnf65ql3407joIEjelXZeDeRHGB0kBV
3B4nfpeURM56FIJ3EvFLXxyMin+FJPo5j6W5qT6wLKqxt8e0gWCjvFvlyxweIb58
HEs6rSXZDlUEIFfwMyTk30kvwuLQ/O8jAA0RlN8lSliEhP3AIhzkLbq1v6r6LPfg
WS0fhJtS2Yhm4enOgwamRSpDmFQ74drS5DqBZOLVJP6mXJhrafwdgho2SLezlydJ
hl1dTB1bNr+C6cJ9vOS4kBiKVOYMDAgeOs80yQarS4Nmt/hzjXIAH5zwyipOc3+l
VpT97HPljBmNpKdVZz5GrkpzuuSXa4TwQctcLaDctdXcAuYgEHhV7plqtc+T+U7Z
+K50//dNooEPmzl7Ht3PRdcc1SS2UXIwzBm+jHkhMKH4eavLLf6bPTDD7g0US8m0
8jmEZuM32GEkmF6zT7JdzKmNsiY3duYI0jvqcmS6IbxRVqrZBOKwVL2WaBtMudm6
93Lq5E+lNPt3ApdjE68iYBEKvnSzHIfR50U6tEN1ABQ12Vce8TvaTOQxs5aIe+NB
plTHzViI5UKTmmdi5IOK2h4uYfyd/e8kITtNHqknRGUIwjb5XTuD3tVXOonLypb6
GCHittufyGX5v8XMltBevqSEhsy+r6suWJjkpt8b5naUraefSYYbH/80gaaoSyuA
Ne2b+Cnfnnh+ashoc/adDvLcWMZgf10AjDae30waidTf6rW9avClmw6vUQrk1u4/
pkQ6iVTZNSN8Cl/uzamauXRZpJ/glKtCCrywpHjERCYilO13WH90qVVqdALOfJSR
wO6MhMi4XbIsTGWzaJdL8uJpPpY6nlD5toemX3pUvam0z99auyDVrA6F+uNRKQSc
FvX228BLYbqpYT4C9+3k/wp/48SPGM7S99rPIWqz1vjdAEBYHN0qFL24bAVBqovi
C6++L0LL7exZ+nZmtUZrWK9IU2rAp/gVydUSnRU6Tvn1c2E4uOSvdqb82jDNazc0
NzPxEDTmNdJ/yOqSYVLlSgr0EMBgoC7Uzd7yD2NYSkXI1mN46KacWx9URXLig/gx
7SekFupK7Yx5wwobfA+LGeBit5B2xUwVL2EUiYitd2woJjL8OTQBbpeojRpxHuVa
iLQ2qLGN1glIK3sAk5yBzwi+s2EL05zqRTbPL7Ck+fd3BkZAjrdZGFs78z6s9t6+
5rS0Db0a09IJYXLjZL0xy2FaeP5Xco7aKDutgUpm9waer+uWOE+GyEYpMR0w7rkQ
1ydw0krKCSnY1A/MRoQd5u3ku3UGWReN9VcCsEJwYfjtHkuE6PdTTEKFNNZOZKR0
zfc5iQPebW3Z7MQeCmE1ELtEVE6LaZj/DTG81M/53avVuA1mdcXXON9mixO1ViWa
g9gT+mbU3FuFwU+l5BmbyrjNtPG6ya+jRNxU9aYO6EmE8/VnPP7J623bh/GAuZhi
UUBMcut0cbxd+dGpWE9Zq/KzafW8CRq5+LyTYKsbd55gu3gs85+qWC/lJzFLhAqG
xO2/yjnNtXnmdP54nvZn4aeiuAs1KTklkIEFCdY/uyCr7KBOWDbvuUA1j21+00bN
OWVCFOikV1JtapbjxtZbkGTvv5aiJ0Iu2TPxeDQl9Q33qLHPfHjUuyG+GANx7XFV
qZhBGzRUR2ai36JNs9pXvgVEJMeS4G86WE7M2rfD4AbsCdjgmOqc2Dq56V8Ym/G6
CXD2s5nq84FBpCIMqnhf+MATXYd1uBdTamoe9on/cPePUBV+XUr74cFuwyYoswpp
cVuTyYPiovTK7yApkqUYstQzhBol0rhkdLYSsZz5D6L0U7LWFlOv5zTE+WfAmsJ1
I0quLezZTd2RvYCwV00c1P+uTLHAdl/o9HAbTigiSP/ceWF1jdfwX4xxy0GcYI/u
2Jk8p6MiSpk2MTOZsPXOf7Jgg1y6B3wKL8M68ZQOXLCy8V6mwQM0E48Tzc5Q42aE
t101q2aBOvNk36eJmzgW7MyZLmfaMrEs3DvejigoSttcMja+oq5GCYkBY87ih2cU
UyL4j8gYZPWcbB5Amji56Kw8RYznUtH/Hzd6IzUTMHm0p2JAuLwRccOi8mmYtono
JcnoBxF93oReD7cMcVKkeNNIuptY8B7AGe5H44dFbaH/UhaiAijQxOZxkCp4RHdu
B2M3alOAB6PxAV2zub03yfuut4LAGjH330Uxczfe/O1njzfFU6EItK0Yd+PVLhU+
Warh6a4XsFn1sTzzu9PvsOZ3RBlkALLeeldCzE6lOC50V/Wvt7ymXQfztuW6R3TM
3JM+fUCfJkA1uZgDzrNxqKTnNPiF8gGFEnGHwnQam/Xwefzr13HONFjtXXFSLeMN
5eaDUvrrBUsjwg2K3LNDnV/VXq1HSYJiXOfyGGnl0SYtH+hucTuaix1KDIZVbCkG
Bt7hz2bYgn1RsohYkqxi9LjOBsjrh/d75gO4OOAWoWmX+GMCRHg+WMvXjonaeRdH
sZfuqgFEcV9owYmLtPqyYkWLBhrmNbxxhyUldM0b5j7Wg+1sVh3A44XSaKWuc90q
p5JGaiE/v4RuZM0hAEfpOt/vFKSMQ7/MAV8lUa/nDjtcX71R+czmqTsUTFsAFzbN
20vJGqZvTOz3V/oryJ5HZALDZvewqfoWbbZL7nQ8luPosisBsefkmPtUieagRsoK
EI6wlThCH69eZHo+jnS+/T62HTX91m1Nfu9Q1kKAnskLuLwmdWO4tfJ4qDD43cGw
E+ZqukuXV8066IQB29yd09ny7kEwF7lLx69pgEaAPKaqbJdf7OGDSex6dTzUr+zO
h1jcLzyoLqef7Y0wzcXcBpWoKUqzomcqMisc2xU/CRcVG7bMYcxzdu+oAbbHp5EG
RaQVSdDV3aHT88xNbiv7BBbHNvRa3cXrUkmT4KEu6e0jrq+2V/EXn7Ifo3On4glH
z01OJhRPckeIEJo070EyUa+YMkZAoFHzB+MYPwD3CFtQOUW1MUj0n0lOerHGEvf6
RIlAncrahq1C1M+vVw4MTXxWGo/TKxX92df3Y7/JNxp9ZWITv2rUf9BLMoPo3th8
XgMBv4iwFZlPmrOMssiCRka4lNT7Uzn2wy5LN9ty9rQgI4YLeii1+bxKWcra331m
S5giXHJ5VujXE1APky0yL2qYWbeMEOMHXplFCq3uMksKdDCSI7n6kpLBzwrkxeGX
gYbIZ/msAAlhhXbMVMhHkB1HGO1JLG/Sa7nvWZBdZ/TQsJp+kxWRcUkCUbmuaS6U
BLfYvGK9PTRfyvaX5Z5X9xX6muSEOJbl1pQ/yG4pdRClZ5NSiWrYNjMKd0xnF48s
0IuMqdMIK+JxYuYEGuvEyqgLCbnLxvanvH22xjOzytSE0MePcDFyJzsgCMYwQplN
r21Z2Qiv04LNm1BfOSUdHc2yPN0yRLocKdn3SagdofyFfFJyDdKNkWPDW01Yxxhl
f38o2v0G+cfnYOvzGTmZBu3uqNhWdYffdhHV8hB9pvC05CL1Q9+LxLxReOAwbRqn
7TWee2jCSwsqbN9m7PjnXqA7KBKVK07IwrR6ZeURqLPXh/Z6AOyOwr64pSh34zXM
6KZSdYSBwlhv1ZyAxfJRxGxODlzbQQ/5z5yRfCdJDc9F/ngh262J/2w5udHhhjqc
2mYo/kkuqTtTMJggF73ZPTufSJK8SA1DKXZNY0+HqdI9hniTZiuLNCfpeYlPb2FD
2ZcMQOFoxEAA/71WLCRTLbnJTHs/ulBvRljyWwsV8bB4YMHWEmiPyTm0DHN03IHM
P+6VdjHsPyWy/GR99HCfkQPukUECbY1Wo0QcHEUK0JW0HANA1XxODqh+CaXEfIYf
wJa1HyKjtOb10PYD/myRENQIqt5f7SNObDgXbe+N5w3ELw7L92eQfn/ags4TAhqb
NSupMEWsanGiMn3quOjM1VpNz50+LN+z5FRnrlzWk9c3UezExXy1ssSPf5aIx91o
St/zE+QW4q123UNs4Rwa8HPzl/RWNmA0vM86yf23NDAV1AQUWhdiO7WhzgAXFf+m
5Mk7nrN4quKw8bzhuJL7jvXBNC1aTjBmbFnmPALXTn1x2rya+VVKljokw+iE8BTZ
N1BgAb6LnFLOTZCZ9tlyJJ9i/dFMzTX1+/GsMV5EIkK0O7Ow12Tkc+qhCWmz3/1V
Eo015IQzOL4G+f1mSPRk+xnJqYUDX0HTtg8ONhBN3VeHw8+KW4V/SyDIPKDb7YlG
XnMCjMmD9bL/87kf+XQH/hlSrS1lb5IdhXVAcM/wgCfnYmD6/fflMk7YvYQGcbhu
RyIOv1KM29rnF+d6CmQ23s2QsUpQ03fomVb7RSdq5XUS1Uji9CAUDNTXZdZ18PWd
yUcnm/Idi/36VbuvfTrrvp0RMwEvn/9iTMjv1M9/A1Pac25A0DTv/Uy9FSHiTeyu
F+UkbM/mUWK+zitu18HrMT5XAYb8spDsARzhZ3Or9TP7h6g8Af1z8pJaJw0uu5Ky
qnX7htjKrNIikWaERVnqLOzPdHEE+eu9VlgQsMLoVL8/4quwqLtxMwt93s3+LccK
O1uHp5+rCCvtCpZkt+3Tlcr2bJVpJHzj+et4d2A5XdqOchVo1Pu0Po+XQhFBQOxz
apWFyNXFiz3DuRZ5hOXxf3yKu2ALjrvV+xio2ZhFBS6xrfpVhMBA1PNhnFxK1AMN
vF1mV8FkZrK9R07J/+rEyJQ9K0GW4ukjO4P23J+LFB7AtHuIPhm8t9bde6Ps+5CN
oyp+wrnhx9+/KqL/epDEpJpw5vc+RtR41IjvDrXPVnmKtuTWB/1/4lCnDBQev0av
jJs2KrlmxYP8lJlBeoJCkrU4N76EJ3Wwm7IJnYaGDLbyA5vmLeeWrlwj3Hfq1g0i
dYjUfYsyk6wfS79Vb9t2CNd6fimgp/jU0yHH0DQ3U41C2NRibbfktmZ6+M8sUMkW
1XQ+e1L4uHs7CHaGPQ/uc3HjokQkNYo1bOd2qb40Qw7NlPPkbl1IyYwBFtQCbwbk
EyFuytu1Rv9AjoaFJmWEWUWOh0tTylVR/K/2C6LLSt0yNIHKDsiozNx4BSM1yURM
fpugL6PhS0Myc2yWZBWADThDxUN5MIPVgRbZptwAcYG17wkB/VTXrX6FIqXyZ82P
Bhs9OLk28kUSemKGakT2IqmGJEwRDAHJvUYhbVfplJCgdJiDhwyCWV2Uq9S2T8PG
cebeDkAJg1Sve1p+93fl8O0+9fuLENJxDmD/CIgO4HDl7y0d4R7o6ElQ6OGIQne3
IvYcf7fXHXgrIlvcBwIIjvgmkqnx55ef341iDmTD607sWBJuHm02mJrfrB2i8ujc
J0nyp9kFaoApfe2+gQ0NZBFel6g03hzo5nlJICSIcciy2L/XfMVuQNv7bsk9dwcG
r2tWPa9Kwo4NElkqiCmzzhGRGbIJZl/wu3qCDLrMoKqdYaXI/z9TcgHEYeGjSn7+
DuJ89jZRk6843K8wQHoy5S2mkCfwrm2JDjgdYLUmB1sO/MTS1elPGvMu/gYCCYWj
oaHd+pd4hC+0lDH/kx3+kApe2bVm+oHVYYk+C5AX4jjnH9tG0frEbmbo8LwLZ4qj
lCuH47yoUcfGKCHFgwHmx9s8dDbKGLcXv4RIShlrXOngXmCuMigojOkmA/icLvqN
NlyNgNx4Tuh89pmazwn1L8aUyrR9cbDaRuz/ai+Nalqkp89zbU37iKTlnO3gE/Nq
+ozOsBB8IXoil89qifVMsU//p9PHzllrfoGFrW7lyqbIu+2PM7JMi2d7pWtM+k8Y
TeACjYErNdQ6C5SpQOtKf6LznAnQcR7O4UiEJyZiLfsbKgQTKiI82WzaEBncVsd2
QP4A01UQMP+aKABlevDZunrFyuC1RIzOSplU31xhJTUoG0E2WMj33YfuEEe130Yn
LgoHZClDs6bkY0IEZtowvS4L3F6NcTjDjwr/w9BwyQTaG6mQa955in1Q/0E88N5t
ao8Oszdbj4CNsY2JLCKVLgF2NxCeu4Kx8eNPUOsF1BHfSX1Hr9kJnC63QlA3Xu2d
84qYpLmD8THPtoEd2b+axmpvW4gBVc+NObCgXGPDrjvdSmOsYWAVyK6k38dFDPes
d/vAB46Nw5XCi6L5ag4O1Fi+/IYd7sf6VGGxJidUMrL0vvb4UPtmJ/V/IlTe6WfR
JtD6oL4Dq5qzdHwQaqqvZ1kiD5hGxNFyZVtraajpcinBaA0W6Eo3Vndwt1pu584C
1a3Hac8/yxNSpTadX7sOXFG8Gld1K2YvEPHLSGNwiw2IAreU2ru3s/2pqdmfuxlu
6C7/DSGbWF86QSeUSn3mTZ/WK9xjqRAEt/s0wwSko4Fy01lt4bx5soVFufk9s7mM
tEJIHLfmXdwB34Z4bGLJgMZcDYTYUqcQsnqZU7YM+oaQgqMAFLUGPYL9FB50ey9W
pYGAlYWRqmWjp//pohNHUGQarnVbF2xIDas8/mGaScToliQ9ewGUWGLDO6xOVlY+
iyzSTyrK4AQ3KUkqAH3PmbNCJDxvOHw21q7smxXtG/p7GVAZEG5Eq0XyzB/Q7BpX
1wh3BZFTXz43TlMgTj/a4uwhP8hyr0O296gyMrLzXM5nFzyfSx5CXm2Oa3eiGij8
H/ppROtETnnwtUE7HTfqgVnVLlbBN+/GtU+dB8QvxO6nW3+afvCxp6i+UPgYBJ/x
orUPtWv9dmlF+rKLi6eNvx5oR4zblWXZ513A8JB7YLp860y8OYY0jWS+aF3a//77
OLDn2d413dRgAJq94keEZEgot6GfLE6gAt/5OH7H9pf5/4uhbp53yqlYQazkgO+z
IkRS1b5/V0U0U1ijQLPksq8XAtT4y/vdfOXu3qK9DzGWhLpyfBoS+PTrljsDpIVj
TUR5OBCBE/bsa3zGLZNetV3BQTmwHKzihwsGdTgWguEXIrAyXPOihmOax9uISF+E
dSPrrJWKEYA5OHcz0Goi6R7s0JU9WZ5+bb3MBmfPLdN/8MzhvSyQfgB+OExcGkcy
1oUBOqp7vsCXU8gl8vXSjLuDmM3MvtAFUncQGjSmxTHLV1DicOsK+wt7/UYeTPrQ
sLBC2HRfSsZYLw2vmOwvbXXeVVh9IqPHNIHyPeCwXprRj4f7SwSRvVa1L6YipZFZ
aLSvx9jyfCw2u6HuLhMKvni3sY8QwhLHyM4pn092N1R9s2knvuk8ZxXkNH9qXrNU
wL8hyzyZfhz3PNMNAs2M1Q3L99x5uQa08JjzFNKzYTMMLdAGe7cO5j9jJvoWur6z
BZA99TjaYXQyUnFWrk226aIucBGN9vqxzzELSgZjAPKHaTABq8IcTGBhckObD9Gm
eV+3M4SUHbURKfSXaXUOBWzXxhiB50HFnAwRMnDFD2o9iIj70rQTPIXB/6sYM6PN
ApdCVUbb/LdYUgonJtdvVCB5oblCK5ehTMuBmGrh5MyI8Wevx9wzFSw3lhhLxq4q
+RCJIetpf3nnsNV3DDnQv8jdR6GR+ahABPyGZCNOMKxIjFMc+8PwYAYXuWLeE3tm
/LAfrCWGCJE4lE85eUcBlG9r+GwPdKEqUU21XdBzVzCT0sW0bw+Cg/7HWXu8Is0b
OLLqhES0kqe/2qHgp74EXqC1UQ1UYTFvJ11mRjZ45Th6HOkjyOGApputv2XEj/xM
JblM7GeFYuvTgyMkyXP8OnFe0FYvATpkD1JjXCwJZru+T6eBVtz6xBlTqqKyARjV
ZO45fOXFi/I8ziBqswKL7ZVWw1rGsXOSA5kllS+8p7t5PVYJcR3vkOkZ7vgGyems
o70oiYKsL/ZLYhIo/+le8FFZBttZyUEA74+lFVravn2znVholNry/XgdJWyFgf4R
toMZl3ZL6p6l4zitgq8X66kCqfoYTk+dueEul8cRooszBW+vEiEX75Fxs2MknQKc
YhT6fBZFHYR4AoN11Mc1kep8i5c2kEoO4trrvaefSEmGwriju+aYqTteF1wIIeLY
oUXBAGyadBblE/mbECwV+wzq0FDzrf3V55EymrhscUzkof9Hd/RerEmH1zfjp6py
6xJs+wRAh9KVdR0gTMduKi26gvTX1k6g0N0x6v//te8NVlI/kh0qPG4xR82Xm8dZ
HRqbpubmJqmZhSf1POi1evoKWQterFTwk9kpDYqAN4vmYpM9YZNsB+J2yET3crPB
1pWFbTgIBO3icJKXzHFBmXtmn5h9wk5R74YYZ+6akNm9r4wXn4x+qeXvaYucsO2b
Yb04qFjXQLQan5a8TjvuXBsRgDAahnPprIDGdMdAds3EG1Poen0WwmJXwTbMSLNc
v9YRuiSDp9BPXKSYeDvZZBFXLc179qrBlUASciW0W1FBD/WarnI5SX4pb3SAxQIp
UQvHbqFArsMZkJ8m0BQJW6cFqU8trFQnQztdSHsW124mv6FAyWRUlS9Zm8k4Ko9T
9Q6WVrvdLHOdQ+u0f38k+Yqk0cIpB5eizvBlHquHvMAshF5wLV2ikGcguzEpGO8p
1IWehLwI0WaP542VK2TqPEdUNRCWmErWK2FFmMH1XcR149Feq5l5q2CPcH0G7baj
LZ10scW05a/dQSToSIc6D688qSqtXZxsZZXT4kO9ah80/ucAR0Jk8swUfZI7hAN8
L0zNHtsOesVvo4eV9ecyMOgxvY6PQz2Gx8GVStqSGcJIJy7cx0c/urA93hdMn2oO
NmcYpuWA7xStKmTYJUHJdv4cZJqATrQMM/jnJr/aCD17+8S/TgRN+vegQYp37ZNp
kWOdbIIDhIUZYIKNQburXIFrYNt6WFdTA6xneHJZbD1GLFM9lA/vNiZ2vQvEU0nU
ixPK0lRgrnMbs163Zu85wrxS7RL1B/cYY+pCvpaLEoQ7mPfFQC5hIJmtPMURNHef
IYK6DU3TAi/ppd4Xi7ZmnRJFivQApGLHrnbtMasayJtoSIhYeXAPZBKbAP/hif1Q
yNkuOIuT6k5cjtGgt2vbJSHweWBk0P+G5BKRqDKm6mp8t/8ekxKZrbvhGz7dbCKu
UFO+uplOZNy78SdqQcbIEvOPtTEVwnXvQqH4yQqb2FkpQvRNX3UdUplaXVd92V+Y
xUqgHrthQaLGfojpySIpQLIw3jh9jc8cevJZCBekuvpexqFL24xJGlhStTBbZQ57
sKr6gboG+66lYL5mA4Ueb1DjHLJlCG1ogP8fjOjhZ49/dH1hqAfB2rYfgZyp43zk
blh8zvp5HU21zHnTyjOCtC+WiS29zLjr4a87yeJA/SGLRTZew4Ri+ZZZj+u6CeZK
0XOAGZcLWjrF/Wu/1T49YhZXZR5iImRWn9c55D8wlt8c8FxwUVuDl6b5pKIC6RXW
QUVRoCn7+0JbaYvKgabwBogGp7NPzNjJ9IRiRWnxloilna+4pF2RXe+CqmmMt6Il
TS+K3b4t48lLO/p6HzNdORC/Hzi8Izh0T6X7e+kWImZz1He9M2nMa1/yUgigomGl
x9PGf/na5gp8tOdRktZb+pbZOj92uI4yX+WMMgA6hpir4LIxWfFFuL+fq9gGCqZA
06SAtymhCP5GVGThd+G3aJ0+RPupgI3r5F4pPeBmmcqm117BJaH+FJ2i3k/BQvZe
23P0WH/ZXsIcUMs0Bsd+OZIkQGlrqgvMrnQEzIVHrAXecxvvhEOjM2cGv6Z9Myay
kzoTM5atmf2H4687wZn14nI05dpNfD8ln11j6wrhhO8EqCjnBT+YRVU5RcEQJDKY
8Pc0MkJqQESjre1EeoJjCmQxRGeJ+gANeY5Aoey+SvnzPlFHsHrBPxTeE1Cy9iNN
LG1ZrvAHfckeWSQaJtyitTuqo9c9DXTdHm6LLSLuLh01hrbiVk/j9kbhw1MO2z3/
jY+uutchzibxd4gjxUwZ7dL+MJzl7f+Jf5dO+gvyyuibKKkrZ1toJzlQ3IXIxMp3
bQ42PVNRn4Kb8Ki42t/EPyMdVYAavypvh3VGQff6osEVO6MsexerEuyE4BMc+2hC
McmajhEyx9XfUVOGXObvj8uVKivMHYGZmIVaeU8iTRuxZAmV6cB8ENnsePuRc1B9
Fj4ixTLdjaxvwcecwnx9eoQ/l6F8i5SkHg5avSv56u7GDLqhuy72lfnY5WwTRtD7
eSko97BekAhq3gffKBRXMQBlP7wXXu9IXPYBwZRiiFHk5y29cuue3HGD0zUMIxxT
lw/UpUlWQ7q7RedzzwlO3Fi4dIzikZRejme/YGstsP3HdTpUBciJbyIlBTIeXLtE
3bR5CJmxO4PWNn55O18GCp80+hNiPMbldm+tuBWB2smLktIHFjULWaCVRao2BdrA
5RfLXKYepv8HT18E8c7oL7GePighrBdoU6KVr/K0sCZn1zm5Id593OmxG7GNEtaC
koJ/G5sRGCgl8owUPD+GHmGfqqA8WeCxDbpO2zW6ehgnTVlQUTNlMcXOHqgbVTNK
siyeufeBFxGMW28sthOAezziJdy/MFj3nfOQ6xt0yk5XhxQksgD6hwUaEeCuVDUb
0um3ttTVtGKF+DWWvgmfg3WfLLA1Jl1r9KCCIqWTFrJr5pZtwPoAhbcfQTlGvIK3
vZmY8cHSSzQE5FHKJsONtI4pBLahwmjlZ/f19q/D1unwObNywTVoFguIaN2xSzH/
oZtebBIOc9YT6iMdsf+x8r52n3MePXRVXP0YE/11gBktKgDdzg42zH3v5JV3l26e
uvSpK724WF5wxvoD1QmGegBWgWM0LXnKnwamICsiYKPw1uN3UTm654nAqyHKPnms
h19wcKsAckKN+F+5yn5y289bVYpZmQu8yGkWqT8fpdkrgJM1KIT6i/MAK25j+hMP
98pEDvr9IBwpqwNAHA7l9aN979TLMNalBLPsqFFBZRbVu+Ljnu0IvcziCF9glyMG
cZtvpxdFNV29X+XhlGuErVf3deRZmxguyp3mmvRVlA1Lz4io15DwpnxiQ6ouwSQg
Nj98Ra570FsmeeKQMqiZCoPhlQJNlsfkeXKyMtFYiMRBJU0c8SYu+AQ65qEj3TmQ
VX2wRZfgtYeQcRGhob771OnFq9ZtraNnwojoNVN1VEYlRfBjRY2JXQQDg/tNQRFC
l5EzDWRDI8TOcIEmeOzMkDrRtO2LI/s5WAnXHIhe3r8eZV7R2ZIcgaYV+Zj/qBcz
0fgzkuqEHeVQDHhl9+3IBFbZt/KrBZCzZTnwsubCjU7KgRiwy2adpWsBr0lcXVKI
uRas4PDbfUpQtVDajYonYxKIO1m9ZLNOajTv3O87b/eIIQSURDS1L5ofdEUJr4zi
d1uWfnqcljTX9lHcoUJjuezYh6qzeTDJ8He8Nm02+pD8MFN9ax2kVTpz0klMfVrE
W9w0sEzUj04clSOt047FrxUIihAPeFQyNn3d+0J5rOzEhfvYD6XUU3RjdAbNaMzg
2xfGy1rwCjqyriZZLx4oeOT2o8rH7zOQHjm1LxlCP5wzmc0Np2XYrhQHRUf/QfS0
073JT9ehL0siz4fYhJg3hASE8JVpG6DTGm+1WLckGyn3y63ouXf8ILay2faWuZxP
sslVJFd0wlRscPaDZ8wPmiuXFO6n+N2w/UPzYnT4kyT6bvMgv7gKLP3IxLgRXnPo
UIxBeo1aP0Ze3Oxr4UtQflhkUg9YKGQ8pnLeZSpA4HRSetilmtK0QcrMoV0W+liD
Qo9ui3L8xKU1+j7i3x3XlVYwNtQpD1a6pBu4i2FsuOVFGXzRVlJJh8R+Zd8e3SGH
qqnSasiqOKotfUXd2fGmOuTtzAGqoZDR9M99L9u4LSwXzpalCVJ2uUNPVU3vdAIq
XHQ6sYzbG3SmK2HDbNP3DWsqYCtUdL8wLpX3Mvuzw/xuDP0pl+PYFkRqGIv9m7iq
vUagM9WIjGLB2G0FvXJ+X/6/eOzu5fLPLouwaTsi00IWw5pUQWEqmKmg5JtciCuK
H1dcd6q5VagpmeqEAuDaAPUFoD2fCtUwhLP/0ljMbKZevy9pqNrYPH/IpGNybl8T
aJTt+EkEnc5gJ2enAYpNQW2dAjC9jR3uM/jXR/sjST5MJYzwMf0dxlWu/cHg266Z
LneJdj6vQsU2FszsDQqooQ6jqggR9pirUYNSW8RYl4IRJZhQZG1Hl2P5HQoOdouw
KEp+qx/PVxdecMXVYH298IFuxDkNBGfMH/7YNw8DSVnoYpk9cNLDmnbgbfAHOQb6
GyMYC1yGAGDzTmFRpWud+hYL+mFt9/hodad4sxpCVEpc/NKqXnwi8zyqHq9RIVZK
CpxF3JW5SyUWuDWSRaPifzUS/Yp+wlAYE5bZMq2kRDqFW5iWbTiKZWHWQIbWBBA3
sxemzxGvsM8SIDSDf96TJMIhmOMe+CD88+mHtixI9hLayZQLL0Xf1Gr+UIE+7zCW
AZ0N2dwlZzTcRJsaxLmOqzLLcZ8AAfz4/9XE6VTvjt9ZM8hfw+6KKHEm/ucXhYH8
FKEB+b31i6GCHI948tX7RhHo/DV3Sr1osxnJdr+M8hclcoy6jasx0o9fllVH7gpO
WrP2DXE/4oggxiE3Clv9SZIZa46ALtuH8VG+Yy3X52dv8gL1/RJFUs+lxPJ63tBo
fCPHekjXRE2/WnZxWT+sZzOTeiG8yLOC6wSskMcI+OElR5ebdBRyAEDdtyN6BFql
QuFcax0Fbf+ptY7Im5ZAH1LNTvwDiOFvy+YA2N7mqMe2p78OnQHLzBjIobbCYWEt
GX4jbIfr3TFLFr6qUf2StMAl8JBbfTbI0JrlotCfOHEYwR5zixDIfwZwkECPRsf5
GMczQxfZXXzsrsbGRU/Li5AuxBZ6yPVNosadTAqQ+L+XmhitMAOl/tueyPlulUxp
NuM6sN6BFwZ18VwZqR5kq+W55/yiNuLzyJ7gMgnYR6/BnlQEo1RSix7kSBwxjVbL
rfi1ScjAc5fgEleGSrM2AaIjmf0fKm2FtyBwBjae1GYkYdZ7IicUQK+aTQRAND3w
MNxzBiXkm273eKqY+3pH5CZGBZzcIrkk1joQrABCtaqMvRhINI5/WmARQ9rifgij
QYgVWo0x6ObshiV93QMCizxykK1w1s/ff/z0zIdnbA24wjnxbhQHRLmnuHzX2A6d
wUqbY7r6ZXmhFTM3jJFUwIsUso7siDau7ZRox/AF4tBuurxPMTulFMsVPOrgSCYm
fDa+IdZCaV9ov15n+kee4E8jhSd0fgNk4ZfrMAHc51ALxXk96sL9HPSZcGdtp3rV
SGGlnYOsZHWNiE7ZN0mXVEOhtFmoSS2qMYplUc0Jufg+xnpM3uBoXxau3dm7jrWZ
NF202Ssn+9uJu1sQuJEENMx14FI3HmX55+XoZ6UtGgafo7d3ribdOXARs8UcOXkh
lNiVSx7JKEGautrlb5uKcBcAtGsGgxr3sjrzf6O2LcsvA429j26z50/EgIbmfXvd
4I51AgbDJHyRfTp+zCemcO9t92RuyMvQff1F/013edAtY+3qFh3zRsO9hTHMvBhT
ftarLzNKfMgktmGHiDiFjQK90aK+v6v8+iwM6COnY4+6jn8BtdyImJ2Y9IMitR50
hbLKrCgJhr4vrIkRK2Qtxz2J+vRw7sV6/9T1TBGydv3VlVCK5JfupzuusuwABTtP
na6DUahrffWqGvKdVFIciSUzovVmCFWU2lVz16yq1ARWnBs7DBVlMNpTafbV6uim
Zls6J1KqyUFCT0uh20hLuHlGBGhiEeOlWl4g+t6cO7RixCPgVKea15Y1mHTNqFrC
g+5NIkKfN0tY5qtxsQWUU+tqlah9QL2ZM65wPAH/D/0EutcA++in6DPXtIooF7f2
VZ16JwU1mQ7kjIt6xlzSsXyJTAqTYqSTO1XjKYeRiLWu/d74lKNKKuJJ2+sYHk2Z
83srddsP7OaRqzNNjvRVFXPhaEq+L0ylE5LhFYyOD47d63dFXH2xHJBde4wqMuke
gzsSxmbIbiVPfQgpbD4p02xSJIZylrPil5LpzrdhH8Qo/zl/AiO8Hcp4e1yu7+M3
5JoQuF5RBwp8McVvQ8m+T5nYrNnxFcl5ymer/EZVlttoidrQTahVnqKqIIAjSFyE
l1qKjF0C6k/uZfkV+GBlMTMUtRe52A3UKmbWO+3Vk4kChkoOe/RMOJzXn4oyYfl7
jvPM/O92J+cs4gCK0THx68ocUr4H9qsUfZ9LYzfRNNstG2gCbcIqpmxdP6YWgzOB
4IT/N7tJdCADNydiW8LQ/CSF2YJ8hDsG05c849MGEwIo1KgJKOof8BmsyO0vxsN7
rUQz7SD9pXv/VfQ+RuAX1OCzaqOQJ3ZeZrRWl8rYuntXeLis874wvr81wbDvfv3Z
93fCMnrU7EebM8hZQ8fYpAozxXH81QDfo6JmDSK6+cppZIjI3F0Ypd6tZTrsuGqz
EVknK7KAmRwfD16HVPQYzKNRW0oY3iQcv2W/EpbkGqF/YW69wfBEcYZODxIJnfjn
UtvS7v20I0JNRngSGwBeYYPkdUCHLl8dGH4a8r5evZEedKlndOnTGjpZEHuc8WwT
/8zLdoWpVA6GplZSkM89e3efK0xrS3pMXVrXO6nbz+NL5a4E7SKhzWsGhSJLDE/V
7NcDt9bb1y1TYHtXFa/Q11r7z5WoSMKMM9M6vydl6w3HIuj+3UtHLvbxtyr2jvKR
auHdTsGbMIGz2o7V9iedvJ0BpJYfAoKnH9N+2Rwx4BAJiWjG+Ueg8X6aNpMHkYi3
nBaeCigxjVElCqr4VZeCl3CXSOIECEDC4D4gjeMU8REV7poq+/p9+nE6eeS5uZf9
51QDnHM/7UYnc8xgsb0jZYnWDkrMY2bJESt/bTuikOCd0/s1GyguoU9AEeqnSGHK
9CaENioL1JsdqiF+E3orcmitmfW6AsB8esDop2NDUUcm8tXCFQAKqUSyZO2+Nmx3
5egnaG5Q8xsydIe2S0h/MeD/779JdIm6t2Gcz8ikVoOMdfPUHAg75SjSCBj/fhEK
ysXZ+4RjjHsl6rWroBd4+p/2T/+FisPGPASlqScMNaLtgSDIE/P1mlkFtDViiU7h
DHNgxzrCYbeeDQoH6zm3xc/7P3UvO/rL4kDI13cl3ED+2Gcmvf7TjRcsp5P2KB7/
J4E7QNbA/jyGbtTo//ZVST3Ef8pOTGI1eZ6/elM+E79ILSiSRKFV8dvDJGgSOuAb
kSX74KlslBe9XeQOz8EStLO+rao5WGrxA91OdycbZZc6qD6qFRepaUHi5UTDFzGQ
kx8bynCMfhIChkor0TZotO2PMZjjO+YbzhnRegd+XiGn57h62/DNdEs3VuTgn/4u
Dvs85WmUFIcS04oMYjGgOp70/iz8loMXhTVc7DNcVJYlvfjToPTbYbE5RFmDPhAC
TiYb39SwYD+Q06Ov4q+KGBBJCxtzTEjyBE+yBKFHAJ4qDVMZALVoz1NA7fU1G70i
KCU8VkvP6v7BwSG+XU8DkQZ8VG8rY59DloQRY84uEVAZkO0pWsphLLSvbyWSa1u5
bYyL9lZv/UIBhyDqP9T7d8xQEMVyd4moOI9hKpUrC2ko/EBuB/NAZPEhNlPG8sbC
IZPQf86zlGgi3WHUwpTw+9s57aTpyHJhqUwgaKA5MpUncwukr6EFWbIXHqUkdwf5
+SOdpMamKEmRySyurV+CIiXXuv9jUDX9l3MXZXBKGoFNx6r56S3ox9mES2dQbakZ
5+H9c9DcZ4ShhgCKUxdh6tIakXrl27yTVft4sERG/u1UmRup1PXEonzfghEIYf8I
9TgjaOA/yBjrFl9Bvst5+JAW5NNdB82ZlLAP9DxO8U0fE3L/UBtaKBr4WFZ8y+M4
iSfCtIc8hKHLAjMFNl+SbQS5XLVzeFhMllnQGLrYwQHRWZZ9GOyvqM1XzJoVowFx
o9Hkd6xc8lny/IBUHOBZTkf7usgAveMywdNtIzhHOIiJPuCzqTVz1dRpn/6C7zUS
+Hh5Qc72W7VHM45S/heOvwB3YpJfHrubXDiOatZNcjg/w9zv+Efi21a0Krpx7OIl
eXdn2J1JfvUWUUziMD5X5NvYe/3jNMoWbJfyh45TDfZa/2k/JdHmqe0BkGbTOpog
WCn7Qbzfhm55+vmA6TQ3iQRnjZpYhU8pEn8Lz3fV338+UNMcbjED60MKJE9Pmq8t
Wd0IWuGFFMjLtYVA6cPisdqb34yAfU+j+kFTQUL3TfHhtcr5m+HwvQ/N6e9p6zwZ
pT2+f/Jn3XayKNpnJzlki4tMf/DfNAdEWjSVq3XcIBVrYLJrupat+YbF21sdGPhp
pSIfGBhp6tcnf/0BTelD7GTBPzaz9nouz3P0eAHY2anBmlZmg89v8fhpx5EA7w4t
uJCuU8RKNa/4uyeg1QKqeW4EiDlMjkXUrVhqnM09fZybU7W7JPiULMNX5geqfzwc
5xJws5KirG/vzO3z9JModH1HwsnW1H3qCksLlstWHdzLcaVJyIqoZ4fOvyt09Xgz
/lvzadkm8X/+SBDubfD1B7jG4qkPNfshSQ4bkvBeKBeBGp+wb/BWL2sHUFqZPqgx
ER46kDsw2qtYbZdBgzPzGwxBIY5UfEOPFIOGfxw6OBdrOzQdcNKbJckzOZ5KMp7V
aH/7xG2JyjNeiiZaUwoA695sCYd27OWxoU4SjBFiPxmW2rBanGG8OiXx9D3Gg0Lr
7FJ9+6uR02ex49cvKAGijz1jQE/peMZed+bKEqLj06wUcDzpPdiMbiFCoa2Mv0XQ
lPNUF0D5i7H8ZM4MucIdtQtm1m80TAX+CBYzkizmaXFD2539Q8k+ppGKiQh5gIUh
FDi/kz4m73uPjwW96Tg52tkiXvuhLgXxWE6yH30JngrAbvRxlMN4n7a7/1N0ENVZ
aGUbTbub0HhHwXWVKGnfOiy0WbLCxhdnN4whGOhF40dQvht6v2vIcslQYFw/PMr3
Fq3IYFK+IvMED3RrdpMlNOqlh9rv1KpwQ0aCgiyW3TBLl1m1PPrYo/TwqNvwsedw
84w32ST3HejMXGNmoOtDroQB+9M1uQyW6uQo7K4k+yAXmNh4VnkY+CBSecBIgdFW
d4fHXo9fbnj3kiKfgAv3Pd/hNmKZj9GXxeh/5+2pHJ/k8G636l6FqVmDoj9Pmkyy
wgp40Gn1GVsa/f6cwvdEgQl9zPUTuIktG2hPilHI1uRXyVEgFQva1PK6PIHGBmVq
AmxWeq177tOaZhZ0yeOra7rC2we3qYZcTHoLRSO076vPJqDtVlKnjgsea0fIPjoT
VC8atZLFzAeWdTivSRFZKzet/HcB8lAY+y1kQpo1wJVWzAovPpPlnuhrkp9N0K6g
4vzZ1k+tTTk1eNrnYFdIfhPyv3TNw1yUKBwOrntM7RA1EHYO2aK1i0TKB71AY1SY
WZVs3paHBCOOH5mqCAGzK/xfXvcY0ef+BwCZoDiW3Vlf+gsCQG5s2QS9S/5U5u6A
6OdxgF1ib6KVy10ksyr+iMHjOlgMH08LReoVByyoc6IL4qy9WKqsOnPvpEPxY5lp
o6zMogbVq3w9mOMH7SQaEK9I/Lt2spajndwCgrNST+4rDpAuyVvOz4gSOlweSqPz
uztrZcGWm54eD7jraAX4YVSU0cPqg32V0tu+//rIVPIljhE51IZHqXxmoYbRAa9v
ZeTQMwbuOVwAbQM3XhoqdMes80JIWj2Bq+ZpjpahL2s47QGqLTL3SVXKE5+XAmko
Frbn+6SCd/O+SCTyWKVKw0lSfsOLWMRNyCtEPQ4qZXUuOOI/3EPXpeNbtVJg2tfS
gYKAxAWYWwuDhydNT2wiesTk+CGP0cCTOCTyDWXjp2U14T2gRduNueYQsXcVY77I
eZt+aSW1J9uuvYq+IqkecZ7TR0dxtkuaEsjYaqTOTqcNVrVug1gdRQIeYYSrMlKY
adiSlkUIhi9IPfCBIsDyoHyNkLEOCp+ikJcUwU6Jfho5zOCFS36pDuh4U6rL8zFC
ybh0ES1nDEmJKTYEwPKhoFVBQw73qGk8GhQb7BfppiWmhg3q2QpYGD9jn8ntER90
apZJK0zcVwu5GGYuOQH6Fmibi+CqQXBy+DHCZf42DkOKKxqilyzyNRWAwgE0/dO1
8Lojv4TIGnIkfglcSp91ls3kLX4uKY7n6pEhnlKFizA9wsXv1wp/6AbSSmy124i6
21IO6PsDkch/EkrC75PgJwtdI9NPBVl66wfY7ndPnqEecox6D6/Jl5KqS2sKFWrp
8RAbpqX+JPTFnaGgZmWT3uBcwG9ACQnieLb8VOP3n/gG8vO5yOAypV7BoPa8QnWy
0+znUnd3q7E7q8Wna9IU5eXvmZy3YYIQEmWjapSUlfMBMl/+ZHw4lIGl0CwxSc+C
sJl0zqO98CsDlour9SDrjFpxCn9VFqZ6HwNLsxSgTRSXEMnylqpYLyoLG9lN4IrJ
BFANxTbEIpgP2kteFDP95WQ/afrAYoGt9TR2MenYYNTEE6nH0e/q2leQgL33nsYm
2fEU+FN2nW5pjxUX3JCzIzJ1JqQYgrPMIw6XzSG7+8/Mw6LQlHmF14ufzoBM3n6x
BpPYGdgXqlknHZttnQ7W8n5QqXeq7dA7mKCKnQVTyAMq2Awf7PjnWTd8IU6rUSpE
K6/rQwMxE0Chxv3MORKdQfGrAzNIIVcv5uzzoSvQi4AdiJU/shSPB9pbUlkauQsN
SiMX08c5nLNeiYE3H/auvY8dz+sza314b91FSPk9BHF6wpsPhMxiAMzv+JIX+VZ/
/B9mEbj4OwT7dsE0Zh6dnSEF5H/rylyVCh4B86CmJN/V2AWAjzWUGK/Ib1p1S+Sk
CcSfqzl+b+UQfvllTzCXCRsGOWPoxJ09rAeZnDTZ9ATviBiCh/0qqUIXPkpVtGf6
oYiaJIiRtXtf1M+7NDvFFgYJsx0YGOixJAv7WS+62GzoXzuHtBWcFg2FZHhrLwuq
TW2KKz+oNXd1War6JQ1mtiyJRkxAFOX9eSF4XcQN09jdu20QuIxhd5ZGu/jAQAVI
zG1c09qix6xFzzsRKuLgJ2fbVBKNFafdU4kkajRnTZd/XMsSpX3sbm6uoG9w2kQS
LV0DR6DFrkqNSM6BtO/aboHm5rfFysgJ2y1S6jtjevb9G53tmRMLinS5WO6cwhss
oBJhwttIOgZqum73S4/zfxpbSyGDW58tdFSrDdwG/wftxWe3KZe19qmXs5NoU2Vw
yGep7e/2Ve1SWi5m+aLW+FptSEmDb0eCOI+txe7L5hN3SQH/tBWHMn5a/tgq1xl+
qobFL738oSrb3IqmodpJRGv2Z6gYRg3STqrIKOmkE19yF1QJ43ER3hnt3/7gYM29
IGYsGj6qXuvjWxPbCXYbJJv/kOYAvDEcX+8u4wgN120KVSV1Mxx4NKf5j/qQVcsF
YVhjlpWUk9vKPI2xUVHxq6u6L3+y52jzfjlncnu1gQFM/REBggQTBBQ05S0qZaHZ
film8wePOkBKc/KHI+2l1Rg8NmHP/iZ7nOHuqmppVDjIYBkvoJIcfN1bRqZ3rXtx
Ob99k2G+MyVPWJ+td/gfmorTxuPZHCF/OzaLyKJE1gn0g2OpSBSk7KdF5D5vGq8S
QpmTzD84IKt8/QRaWbOIDJdh21d183X5EgArAAqqQ/7dkuyBSC4S1xm20eFCixkn
lNLrglp9MrhqlboDBm+b3PeDsFvfjIQzEb2QSThYNjoPO5zql6lSFRgqnfMZ/1jZ
ESwMjOqE3FwLLxH5v5Qq/Nz7TzskKQyfwiDvVULjQ6USU1644/XdSmtaRJOFZt5L
Vy3nWooFVQbulMd8kDpQLviahjroHnMwYP8rRetamRQVorj9Zgf3DvKHL/zU3KEj
ttkKm8+9YAqN4nKlhMBEVFB2/8plce2EBse/2NOPPNEdWdn2Zwoc1UEEXjmh6MLO
ACH5wJtOPg7sAm4snhTTHAwRzH7V2J4WAZqqcLiX8BTYsFLLMi+L0uY2lKi6hE8U
CGiNJAUXztDCn0ALF8RgseZCaCHx1pHSj7/7c/eHj7nnh171fGmtKH/9SS+yLZJM
JCkjJHLywWkdMjUjFZG2vqHc9BbxLljeh0wP4PpuknWRZnnIUkFQvMggeTNgb1+w
Crt96yUUpcO3Jjst9/SUms7ZoqHCtCSDLU+7KbJ0bPAWi5TZ9qQTLw29qqzAKYnR
HZds2cYgn0B6QPDsYZlfTZ5nOOkP2D3M3IqQjmGJ/Ofaq9/xUH3CM/S4M8/Wd8nD
N0Qv9lda7Sn5j2p9fsQ5G/xxEas307ZfKxj93DPKoeK3KptU9G1aEMyO9xDj5xQj
w0QMAv2tQBX5xcVxZ7va3Nz+XVh0lp9sF/NF89lutbNmw02qNK0zrOY1DKPtdhzM
et99CIygGReRfvZEWXUTc9uDeLZXJtQnET/qgtrzmvS4EVsXJS8c2fwazs9UYg8Y
6x7qMVXqLkExROMckmP+iy6Q13lUbpi9ziBZCGfkhflFyThP9Xv6Cd0vLp/nNMb5
Cd4Z77RDm0aJCL8fTz0T2NeKNnEPYSVcQifRUurQmauepWlkMd08AwJZURkAu3y7
i7rj0TeVS5bnTFuxoL36ihrXyd8DFYXUHL0eS3fy1uDlIfqfoOh/N8hG4/cSL/rQ
eUXlBhGw6UUzq4MzWU6cA3LH5yVGTHIYdlAXrsWPkWYXhs8AxbFaJiHY+Z95muvt
o2NJspjml1e27ACrRdIqgdjtRENZZYzIDNuPFgqLebNfOeWdCzvlZkmSKKyNp9Dt
WOMsLrvekJ0V3NNRBjvFmfNohIqBY0VdsqGvkRkMpGr1RlMFpigxVNpWhZVvTpX4
g5scWdNkQE6cw2rjXg4XW2Y3AAgjYxon/ZP0U6YXfP8l2O9d5UEfCuyRYFF9cLt8
rJ1XRv3IrRi6ZOQM9L98JH3SPvUpmUgdNgnZlbqmjsoU3LOyUEAVDzYRWMRlH5p8
MWt/xlivbkWWfrThOsx9XJXmixafkegtVoaySGjQQWUejYPmpWCYif4mmyYxLO/1
aNIdsj9rajBKkFLrcKJ4edWY9/U2yLMGsbwa50zyOnFm9X0YT11GcST44YdR1A0B
SRIp8lkHb5TAsQ1CbyQKqNqNn8zepo2c++iS8v8KmWAAvBT/hE43fyeW8vioaZtb
gr56mZVbH4gXFDEaaymTI9HJ9fSVQqeRSfZhvIgchs5k8Pgf3e33gO6p+N3wdZeG
DxtJtHPIssDtL39R4HKjwf7y75zT+AXk/xiJ9vPnGU4WJWX2nKpOHGrJ9UutfmGQ
YTXx7ddUO3YBM7d0vXvyiZzPpSUPZ10/zz3OmtaB/LEkCBIJPfEFsO6qK7bjqJz9
dLFNMZI6/6gVjOteZMys+qNClots++D60L/PjH++I3YPwDMvQWOGxR9LtAr6Uy7P
5wkBDvsnqQvW5YWXBt2mhNLsx8/2gogbmLKhVi3hVNldd/AbRC9gC+hy6K8NF7dQ
pl3VQtMSYftaMZErMencmaBaOeTKFy/domutc/wkjzIoNvp68Xi0crDDUAob4GSN
e35q6hu6hW8jVdEZJ8xsa6lGyBTGKKPGp9cwkJVeMcGgAxcJ+0TWgQolF7jmaCQa
U11HPxnEW2MgQRIB7uHm9jw+XRjQTf5OLALrj/CkwLQJrcJV1wpvV3bwFV8ML16l
VehrPNqRNTdBuFY3xcsrvSGm1IaeG2P97H1sWLGHCgUlQt/MxuN31tn13n7nxwbo
iY7NyleKIlom9tetkz6Jvm1CalX3EBr1fYSebESBhl31DAGcXU20osaXjRK1ONNJ
fCDlr73+0uGE/yx4/WgKTURwuGa+EcG7DMvkODPAQ8XPyLFJkduYteENVdE3cHCQ
1unKIXTm0Kt+bRog9hpMZB36HGdKHI204+Ma0wneo/K02v8d2O7F4Vva46TjUQUa
1tCPUo/kza+3hCOSJLX/UiIyKnn4/jXuyr8G2r01LzplOkxXRIPdHu5y6gV+qHle
5a5t3+cITk5H3yjdMW5RIybqOVaUYE/uVNpMtX8Am7UDVTG6c3oJr3g6If03qd7h
8rAaACj7I2SJn0WXIageUBYkt2SlEAB1WIwHvDwV5WXkMXZnq45YsCQ6lscCfJxS
1TpHb/RlVu7SKEbCouxRKwXLPnW3ZqFcJfhQtY8p5B3pB0ACXtRTk3J5CQd/40Ln
W62N4njhr9I27uhPOBhalDWSol9qHpIRk101lZF3jiOXSmfSMDPwnBFeV8Noc6zI
TSg39J1L94f0HsVUXWd0Oc8Racimjpgt0Wd8+nH9WejxfjsbfzFLdih2+w1UlUEc
24F2H96gL5XxyfCgfHsoZd4wescM0K39pdR/w2gCPmcANHPET38/8Of5Rtg7tpyY
cYf8ldMq6tZyEBlRCIAKTzUtCh+tdbnLjvC0RH36FxQV6ieNKnoaWVBb8+r2bn9L
Dlf6encIgqvCS4H7v0H2aIaPY5jnuBQMb5OwSyITdSoWPHQrvq1ozeH+Hlcgr0/2
VfnVUc8wsog7ZV3nU6tcVMBfZR6qVRgMUu4n8g5iID0zgr9KUosR2HNf6NJUlW3i
7Jlf67EzT90k3P5uHh2VDDMQpDXFSyWVwJx6B1gbHtn1I2QDW8IxLkinejEJBdoo
URK3taZE2vDm10EQ5wvUvk2yDifmF25EFL/YXEnr6ke2rfW4tw8JpEVpwy10NyW2
dJedoFS1JCut0SSpzxLeedLzGU5rV4jFSdXLrkdCJ08B6bfFw1TzTqWmuafm/q/h
exmQJCa6ziyXEFnvm60D2vfeD02nW5MQdWV4f0qbBKVMwuOU84EV7+8T6Bpbs/Kn
GhudA1p3bAUwDxD83935FWhcfmkn1P5G49UFGjp/KnGC4OB0DvXmW1NhGZfjwXJ/
4Ww02ap4LvrAYCVTd4iRu2B8RVfe3tNMc6HvcFdR1x+n9HxkyIiLiEjUiddilRiT
YM04rvxjCNcr+6v4/TTdeKNnxXVcMyruIOE0/g5dYPrFNjKrvYj5wyPoeRjiPFvk
tJeZVSYdGVNmSt9M36n/jp95XxQ8SrnQem13jLa1UQXxZp+C811y8izFqTP64A7N
4ZMFDGN/G5l63n7e2ZYHKWSaUH8BXshtoSbDb/qdj13K/+SAeWtz61clL+mURb9y
LBWj9h4FIl9I6nlAQZJGKDLSknd0tmojtuEDmvuZskUqXUyQnUs9ez8qISCHv/dX
UIznW4D01ekbiZt3r7WTDLt8iCu6Vsw1S7gQm4z8LTdBb/4zwlen5/UGDBJhx9qY
qx82us4jRFk7M9Qt50UzSSS/gK5CJ06upcPrYPz2+v/tyELdiOJKetWecRk0lj3q
LgeX+ri5Do1xKGD6azMABOi/di3/HKAy7SLFSyUWWAguAgK8TuVDN4KETF813HAc
ghqZpputnnyheHNegPzyOSg9aeRRanYvRYdTXxYo/ADdjka84xg4Fz5/2mosz25k
iys0S3O/xPgFcWIb5HH3CSwGJOndZz2pTTdciwM+ZFTknRCGbb6DLze9yVemQioA
2SWv0XYo56G03hyRBUz/qiYDdLg92MuvUz0P9yEirlcjWbPnxDR4pBNWL6tWZzib
oE+mD9DX9pZnxuG+5u8MSG26K4MHKfNDX4C/suJYLkFGbFH8Z8ySsUCGM0Cxt6Kh
KxvhWpLa/fNtRtkKHxy5ALvLWBLzO7h4Cq2JEVt+/+40O5mTVqy5NMF5rpDV+NJq
RixuJbv5UaXAsAQrYuZtJJJH6FeHRrs1AAnRAeoB/y2syurPUk9nyGewiPC4Aesf
r5a+OkuB/wavxrkxaVDndSEd6w/5jLYc6+3ORYlwGTxzp4zW7rwTeDZ0e2RKp1SA
VCQ/W+ecPPv432l7IHeCJj2I2TddFBjNjZdKvc0fL/Jm4ZsTfwln/9sduXty0MQ/
7A8dP8eA/QoKYw6hDEnudp/pBMoCoXTfgdxBBrJF2vOgKx/iKk4vnYxAsT9UGZJo
V2gLsTqPaPQkEKDTyhhwwcajyR5pYQpyFlDVD6PA9S0UsDk6bvA3ysjQFonloXog
B2ONahAsS+/ZiG2Ah+o28hKJ7Mnc+bOULgUDDhwPr9r9O5m99TfE8p1rJjNuvACI
SiJ3ZGU8JlKek0dp7ifWE6PxpY2/qDivnOsj2SKnk/IndthaJsA3Yvj1W6fPp+Ls
h4siog2V89Di73zPSy1BM46oedTaovBFjzSne1h/b2CpzqG+kUlU2rDFcCnH6CqX
a/og36K1R5I7V+NLLzIAyxbsnhrF8uhp76HNF1sF08hLdKAeRYAmm7G1K+Gmcz9E
+HNgWLVfFUVqxaGsG4qmyA/s0kjr/sFsUPftqcrv9zRaXlxjNrujCFcxpjvJhL5f
O1qrK4Yk57ZDeUM77/nriBraXO/BiBMJJkPjw22NwvES9HBFOpwI6N9mQHhPJwod
Fh71GhSX9U1yXZrzuPUTdSOPoLIcD9aqkrx0fFoA3lbtkah1ih8nRYf6ByxHrHI1
XRstIybDZ0gTdynb/QBz2BkBC/aai6KFJRWH1B9z2quZae0HkZhQSQXr6xwTiO9j
7rD/PhnJ/1jNCpSAPuJTVsESCcfCRg9cnt9FVrUElNBtfMN5JKkBvpfl3mhm/xPA
/0KOAPPO6ZBAfLS9FRGSC825NseG6IumtbMvxd8N9eQHsQDyNhklhbRj0z1E4GUy
bj+IpbGakuIgfYRSggZR1UJSzMejNshPU2ni6aUSz/R6Qj8KbybWWVm6V/FzZq3Y
hlDE0apFvVdr0PYZj0gzC5aV10vqEBxz5LPdg5Y8M3qheKpbBqW8oKPAc5ByUCIs
pZQSm5na3GhSF2c4nBo1PHKtRohCyJTqDatbTahc5g4EO1g0W4n8A8ItfSCJjOSR
i5a9uy2Ar6qnw9DJbFvhyyZv4QbCoW7hi7SeYkgOvY+BcaAQpdGDjQ/wPM2FVyOY
QdajotA0ktddn29u7pT6susxPSFzBo97tTov0jIfhiD8ZIr04ygVEw5zNFnAZB4v
qzD98lmFOKNnquJ7dGHWOB5eoV9g2myJMJ1mmv+/7HifIq+2GWqeNXst7CZynsls
pm9MHLqRMbmUwUuXW69nZfwT0QbmSA23U42Dc8iiRt/XVbr4GVaLXFqCmhyJBJCq
nub3QcSt4EcBZ1aUvtogYTtpp4RDPiBYaBHvSK/L19Z2iVtZ2MgwaklB8q90LRjk
VkvabLwu5em5FK78hymSvF6uMqQ2G0gdQgPeMLY713UihVjVGEeHtwgSN7L1mVnU
M/OHMvDsQQHFWbXVBUDbNLzGActldbl55+ToSWY8lCtkiDjR8+hLUdKp0FLwCyBb
skfDt9cMj9b1TIHkGHr4/VwUJdi1kaWWZY/m7VA2Kl19YG4z1tzfpw7k2hG4OyL4
q7JuXw282YgKkJCWnbEZly3+CuEnMYA+/R+crsaFw46teU46GnHXbU4SDMMe3P41
ASlZxReOZHG9AQCZkL1zgRH3Qt24+vbQI41u5Ftp3VuefNEFRu9iO6StPlNfDhl0
jbHxWuS1451YR0nkORGomIWL/5yvitdKI6iT1ZOSoFW+aeMrc7nuk42rviN6VWJG
xqd9C9iTTyE0kJtvVo/X69sr1U4hS9TvIF8NNcmLqg4NvCe0vA0iTfCQzCrpAWzn
geLcxGFC6nSMpnxUWnxJ4klx0fNtgcJOUzSaFxAgBsfKrXmLzCcy0eU/nWHuul1I
UDPAks5LfHlS9+4q1XowV5nKe+47eJQWiX/Dt31f8SOGUWcWbR3yKszsngYD2JN7
Nq13+P7R/P6CCgB7OIdBqXqyzSYcufoDYDZyp5YtqYhaTpwwpfcwsuNRB3hLiBFv
ypuvAuC7eJcb5eCmVuOVOlUamrkk57vYWueL8fHE8ItK9vevrsZVWt3zXWXrt6Pr
rGPztLH4J8Rm8ej7eEbdQmeA6Uz/k4hYW9WA2gQE/DCNjXIQ3c4lQxesPG7EOiPJ
VKtoe3Hme0tieX1ORnGFu71Ue/9Wed7nCUtJFXX43HlqfjNjUYuUta2ZWoad2Daa
mf09JSNVswJ0vj5fHfoOAaZW/ufvKsxytLhKsmxVLQV7i4JYYAWkBxZeSZBkOMrI
I7IYrpah+o5OUajitqDh0ocW3CDxCeix2FSpC6vTMmbwqdVmUcJyNaMxFdzCMiEH
ZhWEW/3A5ZWFvLYPzgboJtVZMOoUcnGY6/rRzLuKM5M5qkTPCIv2F1n0rFb44JRf
pvWTQOrlg7Enxt02oDluaM7hTKy+J6oQVZXO/KZVU6eRTSyexH43wd09V4g7zwlh
4oLFGlM0uc+1veBifOtFxconk2Usj3DxyN9GfgO7pTXdA/u1tE4ZNwLsiLzaG6Mn
rAQNAs9NGYeuiy6SB73TQdJV4eBmX8jB+ClcHACWneIr3KClH6oAISSurtDGlLkX
lEeNyoYRvO25TUNTy2DG9tSZRKPK44LdnBnfcWwib7i77btSkNy1EBkoK0Eu9sgn
p4dTSP+lU+Ks5bcIyNKftdiFXVYmxOSdpS/ALYNCGIIe4PP6tn6JNDYh/JSIb7BK
mFRQyLDStqxWrc6i4UUXduCG10g1A9tHnu1VrB8dioNXN0ZoWsyVrV9CRITRMS+O
V93SHfYUeMqL0CrmoTt/XnoMOJ/++DgsMBs/iOcehgrTbIFD0HGB8tIQl/0Kh5jH
VbR4s2SWuzI4GOZkloBjaspn4Joc5JYLGG63xYHmNSAXEk/TFdrLxnVcYvXOBfhg
xdrUIKPapL3+vgPwoXGa+WUCM+HsTx7VhrtO0m1j9Q8fYWMbcznStwqWqjU/9M07
wZL/wW2ZlWCXuLZLN2Rsem8xnfJ3ExdRtcgqyuUYbesfid3fmWW2wE8/4meUFb1J
sU3ovM0j3iDj+BEFqZNeoDn37qt8kDOXzewZWUxQMui/D8VbreJxnq66we2WPu7t
eKsquQjIwaBUFLxP31akQ5PTUjQm5gBRJDWTkeY/8yn8ZK/PpWm+wsZ2INEy6Gat
CZqLwQZoLkZj+AnOEw8TMf7gh5kPbbythC/mf3RdBXWnSOXQUwmBic/ZEUOPKeGj
G7YaJyC9uV3HphILAgl9fYn1TS0PpSZHIz9tpw2A42kpC7sV76RywBUbBkfmNed0
99Ee2HQgeG5sfpJ4Jj6jpscvMnQG1QvHANI7CkIyvF4KFfGXhl/WNdhGvNDOZ1wI
gce5G4daf+6/3xVkAM4dybgXa0/IWCxlKxhlQ//M5ylcjUm1u5Gi9lzbn+Gh1V2q
NZeON2Po0V3rFxvhj4m4W61dvKSWtw6i+44TelpxU567KJoXkY3V4W0SxWcBmVqB
zuwSwjdYwGQxIkJw4rEtVnIxsac3Tu+JoL8DUucS0mx246Eb1O+1g9wzCisXaykn
rxTnEYmgA3EMiLFlsYbJRHYZ8nNbmvHaFuxooXg4eISBkhWAM1KLhBPResY/tVLN
7biM3doackU1CWp53QNAsDiyBvgZxaoUF2XZ4qzHCopwdubdnLKYPhLHpv7uOC6a
gSIrhDTJtT9w/rIVJdjwM24Qw9tcJPG6ICo4TfN9t0+8zAqfvaF1VdfftIbZ/vSz
qyR7q/FGsG5nenE8Amca4g3EoJLsrC517Y/xZMYWD8va4aaBsU+G1KaYkVI6gu7p
Yol5usHDhP3bXMnn+atHyd2i2Tvq6rNmWp7iukDHsOBh7WzvJEjRoPfoyVBDTmaY
cT43z9EvJPE6WLILGL4uUSs/RKMTFtRsZ6mFh5t2vbiLxIyIQ2OgMx58Fhis5Q7B
9XYjo/ak3MrrJcyZwW771tB8NuO4bNiqloPMpz+gZo5V75dMwYNH6Cfe1aCQ9BRY
3dCWJCqSWxRUcg2GeriE5Jsa/KPVJUCn9kjEQbQlBd+zDQB3WLH/0/LXOdgiRMZN
DCtkBwPaczCvU3fSjBIHdIWLc6LDqfMiiHX+HElEjlznBveSV6hevwNvXHHnXLqf
SGvDMHn5D+SBQqyguk7eIOTZGaUvgM5wDBVaR7ezubZdgR/Siz0aeC6i2sA//hV9
yhPu1rD1J7fASpONt+ULXWh1y9nUSc7uwMbjDkSTchfahe8kq470DEruAMpo3hrH
UtvqnSLj8UOi7AuNaAY8JLcr5EmIYo2jgcJthmMPzLZIVaApHaS226g4YqYAxBPT
HxgrUC18U+Pijrwmjk46shhi8qwc7FmJdJeINlZN1pIqFLOlgIA2xGLMD73JP6e8
UWzT4ykVgl8wqDg6Lx0Ufc1ZSUXCV+qO0rC6X9gOnRESgaXys0nmmCTRUApVntk1
o2LSFgdSe2tBDYoO+2o+Ds9bed/cC1NC+8LkMucWEenGLVUQdk3abWubOK10JwA3
S2T5pxIK+6AcDPVSoLVAy0/IoVTpshi8qKQYH0oxVdwpWfkEhgJ6JYGLY8JJTHAD
CAEJWXLSNGZsaajGJrJ7lHfiaYImsF/epPXKy2/1dSIOUGwTif9w18L4tVrSuC4e
JDbNRL+NVX5oDUC5UoBRXi7refJHCzfCg5Y1oI5/4va8UOOH0DQUZs1zPBmZPYgx
J2wGwwnIYqXPbFF5XbKz9h/4o4bOQbhDivXCffrvLG+ER+UHncChk+htruAXktFQ
nuAlYL0L2pWrkVQHBBItXKonCh/7hZqtkHNyg7j4OH/CcHnuw/FLJTVXViNtj+QO
xhyipQPGxzyQYlSp8F9Gj1kka4l4MeDNUcbQbAE5X4bjw3dln7giN2v7C2cgA5s+
2+bLrEozSVIdPQDmW4IvEnNg4qkccODcn/ccPTDJAuF9ibOKQQ/Twmgjh7XnLxV4
1zWvxct6GlP0aYPej9rhs6QjV1jMWP+wKptmuUuxldJedvtQfk6wsbrjedm0QxZP
znwYiXldkyfiz9u92Tghc8d85RO7tMB5KR24IVK/x2ohndjKbTZGf+HjTlAl8bvK
tN88Pcm4BeQn24y+fMrjr5H67uVYtV8mn5EUGuwHaG33k4EpO7xScKH6LEYRykkp
DK/o9dQrMK+qcrcHWF8d653DH+Y3skm/DeoqKyCZC2BNXPe2zwa9/8gqPedNkq6o
CGLQ1NEvjWKvVVzBC4C+bDXNaIkiocN5rlIBCkFGEcydd4t+ZadlWlTdWlol504r
9WfvNH0SVgtFUBy1YhgTISj2vRP+lRkRZk2H6/E8v/Z/aAXs0ZQoyhrT5Br2KoH2
2bvZnpgn4TyYZWP36lZFTF+IYnPgY4tgbL4nZCz/aGj91XZk380oQq3zoRFskAK5
0SV0BQsrGcKe1ffsxpBZndyGyirowCWryhBEEgi8VIe27RUFZhLA48XnwhHx+ymK
yUzAVt2XsP/4DZaTQB8Y/r2pU6KAOSsZ5nXg8IQeoS/suC8g87gWQalHLl3sg7Tk
Stei3e6najWDD0m3P4z3d7q/DAvIptJ8kOCikXIHtxNRscaxn09Jfm/fvqys6U+7
iJyEhCKFyHvP/WzM9ci4AGjRa22LnrjTczg0JFQRLL262uOmMBgqUI08WnqEW39+
fngd/lvSFMnwHb1TFAD9MOIUPezQn+AyfZ4y5xSy6VH/QwH/05pSuT1by0rkXb8W
CAlfWiOxnUJdB2/84JEub1dGje/dNY0XPzvQ4hWv8iULjkLP5qXNGQzMAswBCrn5
hrHiLBsJ7GPwyar2Ty6swuR5QjdNx3iJKrlxVSfsYbYKwl9eWPg5d0FO4zX2qMj9
ssZwW5m3gVK/kESKLLwIq/gYx95ZoTydaEx1DPVpT2c/Gcf2wbu8nxMurGlzlDVY
4CnntbaVq4I6rdQ5VfJQt79T8f8afPMjVoQ7N9/W7t2w/WnlIsrAJbuWiDXJAyPf
ScTs/v9MjiyI2RJsKoey3cEUIA5JjVDlhU+U/NueF2L84p7L3Ml/UjQ7Yb3s1TKr
STRCkWHCOuPfyyLrzMF6yTuxyeASWnSxY5tiOQIhc3CgO7HGfzcYq/V0vUbjdCwY
F6m8mMd2i2lmPb8HCqv1UT+8ULkr0FnxHodYZIK3WSXOn7VO1QQoGtZCUmrPxWPS
guKYy0LX6ed+KimdTV/1JMY9mSG3xO+MdGRnMNChsaQCgFAwFN+sn46f3oItBwWv
W8P0DUy7FPa5wfNF3ezccus/lsb5AqdNY0qegEJfLFpZz5WN1V/1Dao8xZ+dPmfy
TFCj1VlrY9cFtwGQeZ3LkbxBae/mf784xIdNZguqmV4Ti6rDbbSldPnfRzcQRpx2
MhQ37UY+SS8pcEosyeepYLjaiUTWnT39lvUeF2/tBReYTWKbhhYzE7WyqUCvOZkZ
WENMfSgDVsqjyQYt1gZQ/cy8Q7di8Zifgsd62s6KhIxt7+Eq6cLhbyvkbJhSEz7S
gh08BqRxNOlYURosHhOXQAwQG0YnZrO7PrTBY/7A+dNhjHaARUZbjNhjTtk4kAcV
nHDmw40lJlL7o9E/lhZQ2nz1lLPAJiB/pGSQEJxjcqxOzLjMwcFIFEe6RKGRorhB
GlPZxeK2AtU22Fgn2Uu3fAIzTwVq6D0gQA1OMujU8bqiDmRzB9OMHjTKGubN3zXF
Owv1PQdq0N2kb60Q5KHQsqeg9ML6LjBO5981YUdddB047R+l4f3IVH0qRhyg9NAX
nkooia4iKc34mWB6UxGc5IYn0alVZFGXCcgwKRsxt1hGTIPasUG7f86v3PvqWQZC
sSEhaXYyngaqheFYz40ffwvMoIz1Z5yxmSt1CDi/3jNpdEFQdRwtlbXxMgTbU7ip
eJWhEWf7+TwCmNYypZGQJvElCg6EUK3xDhRS5vxVMBbYx6Gpl6w6uWWUhHMvBJb8
1AlfrogeLOdtnJIc27+3Pc1Ed6kS644PLgUEFyTws0WCnMMWgEfooD3PonZmCCF4
h53+BU0hWz9v8NHBGN3gPlvAvU6ktV5fJRdtduYtgfUleMOkeXrGecD/GaE24Zfn
KOZgmnvgrcHPrNgH6MLAagQZC3y/2sWreOloymw68M9fBvihRVCV35U4HOYPUSWY
lhBVx2UIP2u81FwhfAxVgzNE4SY10ERqu72zrpxhRiT1HIeTilx0YT1MkvO1RFC7
dnkCoQjjguIdi3kbq2xTuvYg/YwgmVQ9e5wSEyVjX4iT8xBuMs5abhg59QOaWgDz
5u98gBqW/q+DCNFYnlYZFDrSLqe3pkWl7zGQnWsGWrALAwhr/R+0KYWtJDcYt8BT
0E6xWEUZ60vgJvdGKeDCPfGNF+eGYe/CL58IgGFs85lgLMLylmiVvv/tlRipkI4m
6+rfun+SyvpTms6xz8gxriqIx+F/IhKhqgR+Y/FQmBGEVzOLBcZw9pvEov9S0VcJ
hioBYEvVigKUdfx+E0WsltreIm49qFSnCwK1AzkyPwAfqSw5i3lEvIweCjtp7gTs
yZVJFHtaUXMRoQ5M/uuX6a31IpQ0PUFb9XZvg6FNCKGP87aDXjtbaALZzbDu7OTR
wQbU0sOlnEEGdh1JXQD1f8k0SuRmPaKE7F37O7HrmFrnXB25RFVmAyE3m3BJ5yld
J+Ziz4IkqJiMSUeh6AmMfgO5yDyUzt4m2R2uWq/D3f5voyBtBLeNkrj3tXMurZxp
5ONj1WWFnb7Nq0/TtC9TGNRBIPc7rHnDnFjdswpapjW4kJgnRvNnqOBGlO2NuyXB
mV7UpcqV5AiLpNwuJo6F0RJ9VQDVC+PPx7lv6gBvLPOGQwOVKTQr40OA7op2OtSc
dol8YbdOwO23IkrAGDFpeWhVOoVLMvF8UyHh7CEU0BV0LoBswU3LpCk7i7UPUTkp
eq/x9O1Yr7EDwogu+oygFUxta6PEsTINT+d4Bk/z4BTDJZtG3m1g0pn7rI4h0n5R
PlB+siWTiqtR8VwrkE+MQXfn6FA6UPEQPqs4qY+/U4Uw7kv0gNnDdOrOH+1OdGTV
IZv7ZL8Uou9tABWk0M3O2FbdjG9Yy9lCPCosYhlxlHL6hb1a6HeSZwGWSGYwMb+x
/F1bmKTguzcqjt3G2DkDRhEJkTTnAOl8o6b+a7fHt1Wz+JUymHy6z0A8p5QMCwf/
djqlHVMQtL3ALJypu4PsmYgCcMp2O0YyAWJX8i7GVFfT6/5gxOC5eOdZSCtGO0bg
ei1HRUNwaku2X3KroIZGFmOPRUu2CJi3Ou8BzWyqmmPYE8JsAy6eL1oHZEc/HPeq
j/qt/l7FXPw9mSKV0UzkQo4nbyievXnsb3tmNPAG2qcWTUETuuoZ112Mr13Ld1NA
69R4xb1FU9Tp7B89lw4+NqV6yKeZOGADPdA8mZBSrkEsilHff8iaY/T3jOOLDZEj
5lYMkE3HBURS3w6bYAslhCsuo5ZfpRaeQ37ClEVp+rmCIIM1oEm5p08j7KE6parK
aPZaEz1oJx5mcHpuu/deQI8dDdW3BMt+T/JyRZ5KiCrbjMVYuvOJvznIUAQCRaPi
lV2jGlc04dSWmsp4KZJqnprx+xqGN2ygNqvTqZqAlqyAf7EJZe6YAkGniA7b4cIs
OxQ5AVxK6QEc365WzIWlpGKJLT4AaTLWarc42mtiTczSGka0LvNdXuPeinj0eLsE
2j3wIr6Cx68r1p4ITWRa89InIeINqQ2TDKQ2XnaNFp6vaYvW9yXhLkLXs0PlfCSS
BARMaok3Nxd2krlGDe3H22pXg4lJxHMNUQcp+oepcad+Y42AD2u6xDxcL2+lgtni
NQnUKbvThnk/dJBQZVp/edGzb/HcsB3j+hQJCTeBQQk7OKJIt0/JSVr3bEyapE4U
F43bww8EPm5ic8zc4hRDRATiVIaHukJ9t/iLAGBKki0mOgVZN2a/WNnMmBkmtGBh
woIwstG1YOlCWstJG+w8BSdsCRaQ5+oD94ehQn2KFidNmls70CPVZxkkhuSD+8FZ
bRdYwN1q01DaZneusRxPqElFYZhQ4dx6f5LE8jXa4rCgyw9KNCQJhhls7kv90eQT
HvYoamVJSdmeJKkD3Zs/fu2Cuis7m0MVaTByvXxv2zR7AaZEvIP/ITpeqz8bLEoW
t76/B0d8LCn70rmW38aPKyYgp68Iokomv/X7q9BYFh9tRyOyK2bjiNyG1h8fBRkw
6ic3KIFonnlThCzIw4yRCFKbBL+xSJ0I90gFH64e/Hd1Yd0Tu1Z8q3e0CbpgpkcA
AGLdhBNb8xGM1HM8fdqDGX82zS7uTlNpXI1JtH1kFBQt2/wgSUoEM6LFjGKnqsTg
UO9qIFZ0af6i8FzsQYtikxhkXKSvqCOHCvgXwvrCMNd1tvI7jirnT0NzLalntxDj
byWVLXDgkSLnipZoMDDE2sDtIrvw1McxeYwr813Kc2tl64+PWr2sOLHVABViZRMS
oT3Q11R3ZE+V2YIcxk++S+bU6AcrkqPFzQLKUdPVh9vDONBVWpcB5x6V7O7QUHHX
OkU/Z/O5XoYk2rST/QRdSFip0VNtq5U4cBHK7+PKo22PYFwmpl8upKZ0MVuwj6sO
zSR+SuUxErLXwOD9ubCnxS82xSMeV9VJ0RIgXoJQ+2pkMxNzNu+ULZEFLsZyh+Pu
Kzd67omehclWODKOsl47Q97hxGOzmsri1uvrNwYCBjnjYOcOLibWKFyAQYw8T/fr
8Y+PCVVqgS5xpXWi8orldAdtJidrh4ZvfUSIEXUYenFcSlbgvT3HU2EA0sjWe1Nw
v3D8HrnAZzMzd9hFGKKLa1rInXR8agkpG4ephk+d2Ml438zyaHLGwU7tt7EvBBtU
fBhYTl8ORFNliHBg8v8EX8vQ1UaolO/T3JDJ8TA0l6jKyVADFc7o5euWwY7NzEXE
qbrJcZSXFfBCg48csm7NXoUiOQF8SYy2I/x1iKiU7f3nWpZgB2KmQ0brP98c7fZV
SkcRfugt1V7t1n1rWvEtujHfPRCZzKcoAxafMN10lzQnergQjwUE4sp/dSDi/OZq
g1QvwtoG+6HsfpXBgHVEoURZfvDDic5ehUalRtZuy7rh2nhIwJtKn+qx9yT6NMUI
Wv4vToN8bllczvI337pLarUNze0hpQtiMuAt3slRUWvRyIsosulVops9Tt4sU2md
4IDABsOcYsLpnGS6hcUOy+2mtMM1i9M7O4xy03DzKHnc7TBmEt7/GMSobt45oEMd
UsCLm1eADzq94nNr/zMgrPQd8o8hWfW1uJ0bN6SlR7KOMnCKJ/luDkzvjlTAe02o
QJqavVvPbkxXn1SSMx8lxKHwbHEP1PtEbPw6HkS4H6aqdOLpZ8PVwfGR8ihD/7nG
exlUFhoubfn3ri2bkDiHSof2sHvVPad/hor4z36lhX5TOI3/oovXgUkmKWq6IzmG
MFycEG9zV68VmF1z/JySOIM9vZQAfpx2aBOUZTmCQwHxYtB+NwPHsQVtruX+U39n
plpdoJFIP9JFtCwP4NATxC2ip2nguvkUEsABh8l7jvZkDM9VWjmizS2MNDZc0m/5
0izWeNSBDjpzg+QR6R2O1S/MXpTHC/6h6d6/W/Z4zexeCeVB9uq/f19+pBFAVXGf
mtQhc/8pAFOQZ2IpVtt1xgP3rM1pgnb2fCkmYY/XGEHkGr2yFAzXCp4vHcx3WTIJ
aByG9r0RjjGOx34gpoGM2bPBS5qhG0o8sR6g4QcMbPAiKMLX/1N27ZyNkvJmO877
3/Co7G8Fhqmi9GgTeA0VCJNbXi6RkVvIG7X9d3ByJ7ZRpxv+t9u/gqtYdKbDooBG
fTAuGVpf0MlqI3B1Kk4/kIZYLXuSBBoYeLzC3NbYJ6N4YZhpbiVCiMjCKkIsALaY
Bl6ZyYbibmg4gflBXw3yJIf1JsK/glPBAeDtjPUsi9XYDqCRUEMsoHVcopW6LkSK
xAYFrEc+Rh5voV4oZUYdlYLV2/VbJ9YMxOqek6aLPp/u/U1//b13YJjC71kV7u7b
GgYWd6gjFYr+nGG4mwY+JnSd2sMZAm/9ERoQ5sNGkzKG6avUMB61Y1ZnAzi1Hxk5
IufWHZ9rb8pfHXXEz0zbG5zg1xPxjAWXrIxgW1wuWpEmAKLSyp8yFt+L/ru8NO4T
SeIaK/YtIrmayJbHkc1I7PYGI5kwhSFR1ALMc9m5zZ7pNb3r8QgyWbm0f5FouYmV
w++vwO9AJvkJKNRvsLaKbbYAqQaGaQ+3VLWEaWvWPx1s/1vQPmtHRF935lxnBJyl
J8iAhy+0Ky5Ew95Cg0CIyGEuxO0+n6CBlfnj6SWm2Wnk3IXszo3zAQKoQXzFjl4F
2dF0T+xrXm8ipGtqEBicSrxpON5mrDxdSxz/PsfnVtTc+N1ELhDPZUGZ1NcUhjKH
q+g8KzIwpdwKIrxzTigwkFaeVko5gz8A5lcaYJ+hN2MCj+1wqlNQVcK9BIVplq0I
bJ7BgPLk43XNmOyMb84oz43EiN1n9i82sKw6idaCrqq1W1yYnh3lof6x9JidpEHr
LsHTZnNynzre+slbwh330BBRpHxlfUNnEDkjgZ+wEZnLTYjKbc2V1UxjtTjFzpvZ
9WvzBrRFp6mVjfv867c+REzzvr4XlXfiojVMXbyznPuVB2d8sb6pC8LfF4/3VIbK
7eL5BCNb1ss7fuQuL7bxLXmcZ5ePEOlR9gE6LI+n9clWxOPgze30hF7MaYCo1/41
SuDW29TdQiimGDDAz/YHnK2Q4IxFnGeT4K7lQGFi1tQjPHN4ZXiTt2jpLde6NZKb
ae3Uv6VC6TBOtx1NooasPZcNlCfThjWfzjuX6nWLNmzP5rTuJkJmc0sKePxbxhn5
RB8g6y6YsZjgZwfXY7zLitPKLL3vddBmckuMQTA1gHl1NrYSeUbWTCSv4ZmOdpyr
mo2ff9dqcNFZAgN+i/vmwjSh6QXs0AhsY5N3b/7A0FjwM6Q2rQP9h4RNQdgQOJ87
Sxs25CWKn21h38OJaEycyVzka4cBGjyLWoZZj1Q7bQtscNqxF9XH68abur8Wxybm
b3l+3PF2fxw67Y97Y4rxcxJkwJVjiwbhRX7SHsZUE4mD0mMt8WS85bDq4FlWom+O
FXQwcfTcgMV2FEVaYjt/HRB3TeZxLpJhFZFZoktRhySTYJpDX7diVaaje7zArh+C
u2hWYZggva5ddvSut/KrEVnFaKrC7uTwA8WdO916Tw2B3AEKUHxeNxzSd3FsESrr
Ih4xSJduyamPvBV/VIlMgXCuWTXuLUoYTWOAE/74kNbacuJUQjVVqKYOn3XduDq3
n+F+lVJJBhcSWynH8XyaBx2dV/dKNq6I16+gLRttENqcYCA9woFGFG1qbJhENMUh
v7SB82cpGPF/ZeUkUwRrwdscXlqjoUgwioBQmlnBRUywTCzKBKCS9l+W11n5msxf
zQnZdY/ck6HQcSGg37rT4rjSYDfxFeHTEDy3tfn19MwlTQf/YajufbQeox75pIfF
d3SQGTjx3lvPfvcnv4vO30kEjVmZZM5f44DXjvzYlMnj/BwF0X+bwMs/6UzEZgg+
egjdtx6qReS2D+A5ZO4t5Kpr4Sxyrr6GXxiCKRX5N9VrX0mChemhC4/SBZW5rpEg
Y2a0qkmZ0x0kyvGog0uVkr5eFKHrTr9OnOulzO6G24+S6h+xBbH9Mb45FjSrz19R
Bz+X0u4MXt66iVD7kKBgj9GV7v4nbfcwkJH2uTS7BoZJBFmFmF06T2izx2k6dN01
SzHGCbEieW0wTNJ8GctA+c1eWwxPgUXm/0QpKnzauSWswm3CW15Y/i1haaF1aTP4
FnIIb0Sd/+vsYhF1jFrztds+24Q1SQARox8S7QjhRY8Xs32iZILdBEOmTMSAijL/
Jxa9Mh8jUyF1kAGLnXwumT403S6LuoTrwx0p1Ul6Ot0io46zWTNAmvXBsTzlT+V5
E6qGF0UlV5onE9nP40tQhBeEeEoauElQWqhV/bSkP3IMFQ95LivW9t23lPSEIk2n
X/tUqqDMsGYO6Qq9sFYPH9dv8ac9TsXQ6MQ9nPYujxONF7mJLxglFEsbbE89+g6b
GPmlm26HaXUAj3HxBZUSQwF7JGWCtSQmcAWS5Us/vx6eUF6BzcaJLkF7NgPaoQro
CxcSXMysBCh/2Ud1LcpQjIixOBUz7cVXEwhmcHmOI27LHOU4Tt4bpqz5wm4q98fD
y35uU1x63NJ2TJ9RLQLkm4eneU3OU3R4Bmrrr5mcbTYokFwoB5rfKRlsjQc0WmX5
yklrWdFI/blo4qX+iHZGOTfRzZNj39PvgnaRgvYwBAQTdqAGv4UMSDW8wTR5+LGF
Oh0IkYOvF3f7QzyuQekmqQmHcXEC0OyiMLpe0uPoeS+Nfeix6dTgHgy3NITuS8qg
uodDvdG+NZavb8bMuLjXmpBLSgjp5/rFA3t7Fr/m+qjz6Q4LfTR2g2HIkq5gAmZn
B2r7LScfhbMe6RdDsSM8UzNlipaHDewiOi6rOyq6OX0vqhKDPLPhWqHgtyft0Dop
qbx6YIJvrhIEA7aGwSaHqKMcoonPZNof9xpFL3zrOWOcekI2EJhjWkOsOQ6UiCGS
o/vEJf2r+0dEoAURYLq8F0KMV8iJwN9l5QZRGC8BmQ8SjN1DiVnO4aEb1YvGFxdn
xA4fbZow6OSs7N1+rgGtdRp0EA50JRb+ckEqTiw4SP4sgeM18shERr4aViu+gd/x
ZF07gNmzi8+hR0TABiTsN+2VAajG36AAAcy6KeksI3vz0hx0vkWcvZIRKAOzFXPM
cHOB5xNxxp9qB1nLizwTdw1i3i5HaoumJOed0cY0FfdtBtCdoANjt1S9pXzDgq3H
DCrnvO9HU6KmgDJDqIZ4VQxFaek+5ZBsfLLxr0F2mma/pQaqXA8OaDFtXXAadm35
erBJbpbae7SWWCDpcu8DOQtsEoxzpBi4y5fKkaPQvu9nvgQrAUVsZSfJxgnpyOdx
g4em37aERgTjiiS6pQ45CVdgikOQ0csXQRdPDcAjC5SnXVzAXzuQaNPe+aUNLfqq
PQqak+HM+ae0+YWeMVYS/5GSagXfxz/FfIfW0Cu1b+NkBNPIfYLIzuIlPJCxoGZh
0TrQNg1qXBgvE5IFg8ip3ZyDKEpQmkg5nEXJLuGUtWGuz095PeK1Z/wwiiJ3lGIf
23zbItCuO8sd0CoOylfnNpB2bluzga+rUypb4Pq6JgB6eE6uBrQsm5XRiI0Uo+RE
sbkmRh0vFe3Gu+2fU8Y9vXM/owHD2OJl7t+I9ESoo0tIyAIN0vX2f9byKz6WQujm
QU7XxoxlngXw0khf/GFvuKu6ch41SDY3c1Fr650A+27ZYGPgmJZl9gaxaFaQpAEx
eAUmb8+IJXwPDj4rYncLG9CbYl4mg71KIkq8GfLan/Nx+oWb8/91od0xFfBmRnhJ
YqfB3d2JcwQ4t5RNHtBjrYgpkdPJfIAXVjRoFZ7oK6cQjeNOxBsOABOME0+Sypqi
Pg8TzaRBVlK0/LK/TkaXectKMe3A+brd4w0bYTZ9fQiVEsMAWLpwHNusFGTf24El
T+guLTlmBdCySycPV/62rGwyhBKa2jBQMJzVXlf0ngHXE66mo/as4iEiucbDlA0x
Ix6RO7++dLY9AT552j6avSux3zopGA7Piccs+Lw3riBP78QBHgnCEwUSLdBcxIS0
UHnYctlSMsrp9WSi7JcyOXiFr0WJvD+1XLLCfK+Ot1cnM85/7ggEtIWqEN1IlqFz
VSxWzRpsqPdDYRslsqAIPPAJn2vOtdItYzow1UxuAnf09r01maEgBd8x6NqDBXt8
lvQoAPEvculNo/xhDyp+bYqR9krC68VpMUhiyay7M1qF9S7fvfvwHhWMPHqL77Mx
hWCnCZ9vGlCPviDA63tFNJeFzlPGBde8Qu2PudWGOgq/K6NZLB2uIIkeiejH0hlX
xyKh/82jmzHPIRS6pAWvjKf7bd+RB8y1QmKgpW2SmzelMORYpjH++qDOTKvrmgFw
L46+WsLsevkwYmVXaLteEWn307tBx9w76AKmNnAFCowolGV2TE52toPI5s20Izqy
II1i6sjl3/IV9C598o55o7K0QwAFgYSBf/Os+fw3pgomQ772B+PqTBhx6dU3nEl8
w56brJPfYVNTG9cDE4ZMsQ8+2M2/Un3scabUI02+rnH/aA5WN7qMI5bz3txPWBve
6sfD7X515A77tN9NoXagMJKhgD5By6cxWaHx6pcRyUuZe1xz0kHIV8rXXctYqAWi
n0U6bNTPWmLkDB87xLA05DEmQO7nCyieooNMu87e0O8vLHeiP4CuZPtPlq7JWIyv
GSZmqFbsctVXk3a3Kd8Q1Z68qIRM8AYFEgQwaz7utAxwrATA7FtprpGu7dcrSI/p
KCnLadfOvBFZHS9xuMnxEvtdDEEMP4FZvPqLPG4KfLiV29CTo0MLXnFFbdshHgvo
+Q5S+QWtvUq5AbCxnMXaRKKeX3DffwKo+OuSSgA0cMlOiIiTOou1vESJGTf5PdNn
gYZjOLB67f/e07EThYn/vE0m76fijQfoK1olut/kFZMdzQD3PK7pkS/Im9NeNoH+
3mREuf0ovWjnRTVf//3etBMVtnB58evQ6toDOrcLyIGe67mh8lMW92vN94+wGq+d
u9tCPG/LhSAlkUksRNVT7ToAnfzCEgW3QhsmJQqALOmmEg9Qcv5kfD1kCdDU3Pd0
GB95Cai/Vns1psBVIDTMyCqoWYPOK0yU6ExJsFRWFNf+Coku6N/akZRP+8LCsADA
xSbPt0G/s+etW/aSZshjVb9PdFol9GG9lQ6DKMdIf6TKoeobrJwr4F0LHBjLSj8D
kkKKHsWWzs76XzmH9LUvSS3O57ZX4YAgACs85K+Ai15DBdlLu1KY5oS/XDsWF178
VHMvff46WEfTae8wTmyVnPM39fWiwhARopx7XJ3PONn/CZSRv5pXUST0FWQtNyb2
aZWes9LKJgdQHyFgKz7ATGG+N0QFRAaN/mX1q/QcuI2BFi9TpaylETHxW+qjCH01
vkaAy/q+4D3X+gEg1aIqy1QCO5sZEArnh9eK3enaDyo/0yhpvup+aB5R4p0uedgI
92vlTu5tWfH4t3vef8JMLzxzI6zsN4UClZLowYc7k74997l9M8pjqRVNndUGuXh/
NXfaDXLiY27ndAlhiVeqsvDodMcT/yrpPnfbJo2OBvrKWu1IDo3SUPaDQggMMef7
mYW+NA0A3LGO36yKmOCVo96AN8LI04Gnuv5UXeS9vDdPH3ODmwW34zxFJXMT8IK2
OZ/Dkdp9oK0R9eb4EU2Hv1L2MFjukBoT3Okux4JEcXM/X4OnG26py0D0BWf2uWBe
FE4E/zcLMvYm4oELjAPHniLO5BSB3jHO+mQ9p1Eonjkwatx10zFEwuWjwguBfNTO
5WcBGSUoWNQ7r3XNar5WnRtAPV4ff49yTmcNt2oDVNMXxU+61SzDILBNgaiYoQ4W
stB9Nr9h5D+meHDvfu+4yF49JVUrCScSO0lPRDIXaBLE+TbZcZZbmbG/GUPvxZkT
dedMBykmJjY3hsmN0LAb47nOaBd9ACGEFDPl1LCbSxhJ+wET3dxN/Wy1gJU5VdzN
qicPkSxYJRQ8mvRC2TqA+RRdyQA/NDrT0NeTv0+CwgJtsvokZboDEfk64DD/MdQA
+SmDqXMzkNtsFloOL0PBKszntJ9CZYGYI4OZvIVtSArcRGH5gdc9jLGRk6mToSv+
uCotQauI/0NZGlWhp70Y57JiMdoWHoAoQ7hlh+88SdkNPepvW4INi2pvbTDoPDz6
3SrSYjkztC/mQ0ePnI0ZJa3/xqAFGEH+psSUY44mEQXeNdefkAi8TSK5OL5Qjg1n
dlEMEXVJhPPQIfqedNvkB77nVuXDk/pqiO26ejovXd8AJx/xFbuUMrqZ9n9DKcNL
OWf884EDkVj2kNeGO0OfYRvNSNyjbRw8LQQYtseftfdd5EPaX//3XeJuxtcLfWBC
rCIWFN3AOQ2wayJqZtcU890UQvfsF4ca+W5wCw8eUSt1K1QGrkYLKpg0lUGXhVAL
C1LSzWJLzkUkRpIUyQYhC/w5KGhxNbXgvQtFXN4d+4M42g4kboIx9sbZoo18cEc6
PxBRgrBX0bOpMptdTgDKD8I/VuvZl1rhojdjbGCu3Xn3C67Q7YVp58/PoXbhP06B
Le1S8tcmcq1ytyIypcVXS0ZkyY84BqHAe/56UutvEgbDGMnDp8YEvWBumX08wMSz
g06QA1xvLA9y2Ho6s7fP6qggSvKwDPqLcf6SPLuaEOElSiEsSdTXTNSwoI7rAWQs
as/9uPRCejoZGvHOKgi43vSpQlcqgjDRlW2xc/s+ptKcsvsVhqIRVrk0sXUTfSHU
ZPvlpEvqMR7FkyolFDexQn6rpWZQggTWfFhYR1axK7N01lQ0AacM3JXADSBKas5D
J7f77MTgV5hYqYJG4oL5C9W1OgHsxiZRrOBPu03uE684rLaBhIOS0JVGeatDQjAV
tdaXhjKGke4jNYWIwt41dQPvi908Uq8zZO8xQziOmLZx9qIcgWVuJRkzFc4XfaVu
EQ234LjrbgXV/TbXcLB9pepGDem+rRbT+svRF7RHd2sErnEM05YNzVtqdQLitmvl
ZdtTZRtLnXWuJpfdHqt/sDT9t5AOufd3DpHUa+czdN+vixm8yP+ZaKadYrOi821L
IR8xzs6ZMNlmfVIMJDOYz2SkU68CcKPC8tCIjdDM6579XpEmPQb0B7NALPxAHeGV
/bdJP1Q/oI/zRXOu9EwzpkIlZF7cXk1UDYcByn8D0dGfh52Qra5Yketoh0EESAPi
PFCP3MrM2C6mCH3COeHirBfAEaxZgydVyoFxvnXpY46If9gkvNxP2FEpWdeTSZwO
vnj6oKS/pFrE/zpo8z+sYNS83ghSAcUEu2KrA8tBkJ4It/ijsDhuGfGMEeVyHt6v
0majc7u60hZDrdECBjz/PjoeAFAw8SpGLxm/pH0//+XsrEPBUBoqErxP1eU4foh6
r7fdTQeOEe05pLqbRxFZmnfozWGn1WZEQbWEgc7N+3OylyhxMdtcx/tjft1PvHD2
YAlA/xDZxBCwlHdgAWYaV2UV79i1vW2xPhUV3H3txeWmxdJaxgOrSEGUt6nw1AgG
hZP51UIwi3kQ4DNZrvrTOh4vBZW/aJA4BS1NbSQRT2Rsx9Cviadp/yZo9WcBfc3b
tJWCWItB7iBfTaFFH9E/EsMR4RfluSps/ZAVT3QP09wugowoEsOqevvL2KYC3Bjq
YvxpAo+3cj1huSFIIwHwFVq0cG5xWNOSouUEiuj1DPCkKg/9tl0IlkG92g4JfxsI
c5kB9jy44Kabu3mibifh6SYFzrziNriuhlFdwwyEnlNZHuW6XU3deWFnpgJhVMqw
449opmJEtpZQ01bzHrXbN2IPd6FQi+5nz5MW8vb4u8Wqx9XnfYgZ2y+8VCBZIitI
NupjiS7SudPmebhsHpXogTouNF/VoUrrw38qubCWlB+nkLifNtWCtWBfffSRzm/I
csK824W3o8fZAP4ClcDASvVRCPtoZkbUZcnR4apDc0z96b4pXtjHwN/zGpkXZJTj
Onpx4Pst9X6+OjsRthdpterjjDvsuq/aU0eOafVd7cBS7vcQ01pOza6lQd/qWFQr
WVB5I0KB/aCAsA7CLoL7qCf9Ewg3901H7opypZRlmu1/+M2+Juti1gS/Rjy4ay6n
wzjKJ+ujZQTgZ/uWi8ezONRKXiSaMxIGiWZFwRrgy/4Xht81XecrEa3vPJFYaAmy
F23yTd8jwQ+NiZxLwHKHs3KD/yvqAD51viK+DGp0ZO/HxeGIB9+1AUwTdtVfkRrf
ien9FfmU50sqAZvL4rOojumiNQ4Sd+97/Jbcaze0Ak/Gw+qMtjBLepsdeZ/oXmA6
tT9IeBtz8/BOaA5svAsqzjJGlYlQtQnVTCERBPVHnKY2O8bL3THZMox+j6GxZRvu
pLb1L3iLZqVW5dAOHX/2MnIDXc1lTvwudgrV2GMhQ9iws9HFgmxRO1AHa1X+/xOZ
lUceGFcarxR7oHyhx6XRQnZxzsLHRkSBDh2H6W3PmNN0k2N5/qjB0yy9HOz8F43q
LYNtRX+46ZPCc1cgC73iDGFlpQZ9lnD9ZGtTaYQh0g958ZCnxQvRp056VcrBf3u3
fOh3dVKDZ070qkWHXgDiJ1FJtcFpm2ia8KSMudp44XWf+MBMvCvoZxEQNZSt6IZB
5Py1fOXzMxz32enEBeInb3R3WsfJCr/LZMP83+KihdpiCHytGkmmw7i4USYwBKrD
Fr3+iIYx6pPSvvkgH1Vp7hwkte7inH+H1hnII6Ino0BwmKxAWGhq3JM3xCwhea8x
RHmSi+CSWD0LpGuIYLciTLARDI/n2pB0v4g8LVI4UNEwx157wd2hEX/wAPwCj4nU
GjSgzNFIMxhlXtmTfOlRRSEW6ilmi4F4vJNqvoHtwYU+7f51u2blGcvkOFoxXOts
mS+vOhxinVODTBapZfK/uqdslbaXCWxUNJk710Jmgh4+zevD55TJdmW3KJ+WHJZc
qRZNHtysTlsQHH7V82xbycPrf0Apur4WIn4lp+bONeNhJKTqvWZxgq2E1nnNskIC
3yxw+vhJT9OHN5RTMssXJHptbVrW6wvHU/enZQdio4daVE62jLsl6c33rD3qyoiV
YDxTq7fsq9scl1gfNLnd0kKZgkjbNDda0Zh/MOdt6DHas6AFLDzCotCALQx73YEa
B9Rp25fpdhPbagELnXf/4iK5aWQYuemFubYOE5AK6humd72E+/Is30Qdnd80fb++
9eagVUc1/E6Ub4Hu3zv5xQ26QsU48DrHUKbZ7F+sQZpVcZmYwUFlHQgD60plMFpV
NkKHO8HmKSEpqzvwyLXEWnrNSZLFxH/vFmSOd8gAYrZ07akRq6ePLRGaifpULpQl
weYbhZZ5Kq06J730wATPbZqJ/nv/2SHo/WHlccaTzRfynJnGJ1fPNMulXgh0c2nz
Ngnc6jc96cvtn0Rf5I26J2XPCNV6L60q+dxM+B79Rh4Rg0+n6GBCapq5XhbK/HCx
+nidx/q9ykGJoqX5rN1bgdSz70UxxTiysddAywDFxZQAU3A31bfYttguqhoDUe5B
C6eROLy50LWOc8H66IoZlU9//c0fowfjJl2a1r0Oetqx+jHHgv1m71PZO4XWwryy
qVxhHKVXOLfoyUDH5l/WGp8cr/svvmZKpqOO6Dl711PodmByQ0TZP8AOnj914Jzb
sXxlHpml5JpbglMxqJGz8HgDKPbGmMn64ELagXeVGHVgnEdGy+ldfZQjHEGtklXZ
BcTPxe3ccZItnA4LdRvZ2pywhegYTD10T42WGiNGrkE5pm/u/NYU3HPkvXJbHhfg
gNmOIiHPVwMit3OCDN6HIbTvPwUjittGghxVydpyHLpwTM921jxRirpOXqhWCuAJ
SYx7nd/oLT3/WNv7BsQ0/aFqfebC4uLoHTXy5s6n/MRSgeQNscpJ805ariiauQUb
NJEzl5NBawwfFqnqkqA6NzWRGn/du8KWSASYuy0Cp9XRCNnXGxiXwIWPlOKb2M2u
hI5K5X4s8zd4s2MCgCf/qgSEcTGNrwxnHJToBnraZU5ROuu4KURNkHUY9se39ckb
s6pjKwZpsM+J2pcttg2xhSfKOtN6Hi5MoFL3fEam/axwQjG/R8u+gRGWpEqWN/pa
GyDc9zAI662lcBgmxrG6n6tn1wTLJfzQi9j1PTKSdMPQWP3f+W/9gE3j9QViqAGL
yWmKmHFWW6XDf4n/y7uic5cFtW4fwlVLQftseNIh60dgzxvvxRby2PZDVHitEEOr
rs88CTEmxRVhJqS9SMAp2r4+PLANaXPV5ZNN1T1ckj2Ss17yOTfZm7bV/f82mwIP
+LAlAZunVTgD1rAHxpafVspUI4DexCOUaxZvz93U7FxgX2VF+OvkKtU/dXKbR3Zv
yP+K6MfwBZydrh1b6ipDuNn3GcPc2n13b5twpQlVmkRNXo+H6noBa1I1rX7AjeDF
RrL2mypnVE9PZwh756MKO1G4ceSaVvPbeSQZVIL1/ZiosA84O15OSz6y76u7GGuz
+Yuvl4P2WKgYzzJrwVMe4cHJBdUKrbECn08azWJnrLnYPhm/Ly+g8wyYIWAX268b
TxD2YoFd9DU6O9GJZKbPYXI9iV7nIZqJGoK1Ym0wzFuF1Dc0CcXbTqqMqJZCnsKH
2nkZtASoBGERLQf8dX11rFMgXghnj/ip+oZ5z+5HSWGO+rgf88HObcSMJ7Svuk4T
GIRe6o9AZVxxKlkxlFgcdL8ezPG0TLc4B4I0ahrQYBohtUxsMoey2crTUsC9c+ZT
79SwmBMi7RMHGhYXut/SN3pDkQg9i53NywT4/eIIWXR4gr7Db7Uzn17e4tpJ+GeR
Ne1o3Z2z6fIyxo9D+Y9trsn4qzST5NQvqz4EhAn5HqNIz8FpMzdESpETqR2EFw1r
BOwPkucjWPhiCbe6db2xvdhWp3HajhuHtmd7XWv66vCxLnFIlzKqfRUnHNLoI1+N
haSEKkhxlrsNOtofFIFVCUyj9ky78hBRW8kz/VAknvXO3AG2PEVGD3hBEdE7qkvF
TKD8RVGfp68uFe5BqRtwYhM7azIpxae4sZCc2FujGdIWRrpUMJa2L6nzzf+q8Diw
TNQO1CP5xcQJ+WNEt7psNAOMkZGENvkagKQx3WwZadJYmVxlxNSaLkfpcoOmttGl
6peq2k/i5mxPENtRVyZN/dGJl9iqlTQ57kHjH+P+MV5ndb8KlCOeF9vvffbTZT/C
4iYCDrJE7pUkyunpj47nPQaXxMvSIMunQfcWidCl1+OKxcSEtwVmWZGGEY0oqFHO
9nCZBqyBOQJCPHlQNbUmPaOev3DYqq39iNb1wTlWpw7nQl1RGMQDRQ/2dhFCEzCy
xt91i9Lzfj0nTKBAR9L7tbhJlHUJHbZ0QS6K811Y8EpR4oMGbcAfBKRyqkdz6BYp
4gRlzHRGH7k08wjAetw0iDsjQyDfwJVCOPiaZM5CoT/BsopRyTx23pEF9Ll8c7QU
jnyH6C1ItOLUQOnWMVnhzbtT7Th7GZyq7hBaMlMyHMHKYYjLr4kf0G0i6MEdHZ0V
KDS0JpFZBHcKempDe3f8EDirS75VRprP5R2tp9enO9otn9gnj011Y8JfULk9JWNY
UVyod20jNYJr5vcM4RfMrDLKYPwARMuyW7vtNvaX9VNPn0mLcoOiDiixyYT5qKKJ
81NH43NHC7rAuzea2/Lse/UyJyy0v8ogg2ilY+CleXGZbQmiDPEGY0P9cw2e7Wh1
ebq3zB3wVGyfUCVnjh/4e8CvCNxyepu8cm6P1UchbIKpYfVWZf5P9ClXXgpZ/ks+
egTF+GXsLnYW6fzp+pJsSX1P7Dk7acjy3G+yu38sBGisniUaYVy/w7PQj6nHkuR0
w+Z7Tpa4hJXpXgS0AiUptyud0e2q8uW9taobOuAzibcIJdA5iL55LhqU1onlIZ3g
+OAuffmrSUhzINd4AN0SixtQSIDLJ1ZQZq32C0fJ/Tk/336poLbqs6JgpwHUt0OU
TmOtx5VWQtTOsl1q/Z3pqC1chjUfo9CD42l0FDCSb3C2UshYWM8Hv4Vj5IDnz198
WjxlMFSPx+/c5lgvC2/biaDNdzw9SBT15BQP5oQugjtIbPcdwnFUuW9pZbvdiCB0
Jl3Ajpmua3vQqSP3HsIpEbLgN2HY4Vk2Yqa2R3kBEIkEMeXlebYgMtwzovBi8PDk
yOUYKk7SYXFgzKSsWkQOAY/SmLODd52blVAjmy1Yk/Hij0jhARI3yq8gJDbzhcX/
joHRQLojoTcE6vxJD/f/zQl3ka3fcaFqZGz70xKl8zj4l1LYhLVwO3+YJL+JcEFG
ys2hK9qNIwHf3bQ7y7UuZ0854MigjVaLdO+v5+3I9xHft3ctvjVQah41/NB5iGOD
fapXSTquhf4hWDSVOugH8GXX4DdyuTnIZxcvU/a4+TvhMoh/7KuS8rGqUaiR6e2d
Dyy6W4UWksrD9TTFtRT2L/3ekfQRl7y14FYA/e7CPX65N3t1VbUjE/irDpRSIa63
nuH9SyY3ZjXiBBiBTbkGhJPIx6c+uQUBlyNBuBue/wTlR/eOY7JQT79Aa+Tq3Z8D
6bGnwgGX8wZMaO2dzWxGy0J3Scd13uwyMK2jzHV2Pq6z8uHF7/a9pVBpwq/UlpIW
OU+CMCLKx0EL3uWOYQQslYf4Pvdo5KULN9xtKHlS+jPbtmdwaqGJiM9P8ttwEwTy
vYMSKgM62MfpH1FKc4MOy6tuWCg8ptFLWHHdPt6BeGGT5Yn0KO6V2y3pRf7ZDQNF
+bXozxqny/O/s4GUnq0axE1z39tLwq/AyNemgVtrXfmy4SOk5uUi0qJ8LtnX/K2h
onx78FhC9NfkO9nwLWQEL1jR9lBnQUZmBOu1mOn9nH8nrvnQWSP5+d703QW2NhpP
4d17iQWrg0q2LvjpCUMywsDd/AXoCPxMm6JirZA5DzCy6pZjmARRqbrd/odCnlHJ
3xCAbZE301hk9c3gXBojPMcLoxAZ1grNXvLPJe1S//s1MWQltPBFmexrX2Tqw6R5
eV+cP2A0lEoBUEdnVgYMR0cem6l6/g5C1IZ6flG+9HbYcWl4evCd+5BwO4aUSJgr
1inJg2bqxRe9D8iNFvqFM9bNKnQ1srWJHqFgAqXlyL1krWbG2YtVPTb0BrRBY/tI
2iJNij+M4jLvMlcuji9Huy0saWCrlskOeCzRy0T+an1ll1tEiDWvgR2DWjfHeHsT
VOOPNDTQ9xqzNX+7nXgNRni6rmVrg3CjWixpQhdItIfoXF+6Dc5xFYcNMr3QwwMZ
EtJ6odJsilxdu0pZz96iS3rIAGZxx8NavlLzOjV2MoUi/AHRZkaf7OsZNaX4gKtV
mDoEPPZQXrefHLcpxLnc1dxu01/C5olWSWKoJkiULb1JvawpfbhnTK5X1uj7HPgX
haCsHyyEaKv3ZxrYP+KMIpMHOgM3rBcQwlIGL9YmEJH6ljHZ2XjETflIjRkjh/Om
pjjECfgdsMtv1o45jxXpK2LYqEFtQEsPBz4qunUICJfr731SHdb7/0OwMjx/oCX3
ylfhHDYDPIr0+08kU786ISWX1RfXfyTxGuzsVnsxl5hbf5QIncDzsWuSe6qm99jC
vjV5JF4GU3IoTVOqzHZ+lPCCMVflXIXhTMqMRxtBohLJH6O1dsSstwmZXEosT9Sn
3vs8RzjfiiYPIqfdOGDvvGWs4mGYPUDoEOpQfE0r+PEs1dPJXAOVdVeenqPoaW+X
8Beb9EE1jTfnsyRbRW+L8v7otfmIlYn1rBmsQ2e++XWErEZLbdiTi1pEl1AtkHwE
2lNkLw4uG+TWXtBGhwBERu6kqpTLc55DiNCkqAnCGZ4306VbCZFbpv1vZ0TH5QkG
yRXR17PKiF8mW4VTT6RHhOETSGpIJFVMllhQC1w4q26SC2dCQ7k3IsoqzySHQW7H
yLZeh5C11sDqe7vNylgFvxhDzHBV0yOrovjebSHjsJXVN4AAkq5ki7ySDW7HJMZ7
06HWXx7oI11dindWow9RAr6Lrz9BpR5EMVfQu7L6WZ0/kOB/9Z+nC0rzu/WF5+zY
PKcflt5+zjnNU4ELjYGvQD29HR62iRp0YzxbznuT9GRAGWTqWOO/ujUWgFkz/OfE
sBlnPv5BwSF0b3TCB4IH/KiKgzrbXEu2VdHXrmnYCrb71Coi7XcWPUHfUuILj78P
grbrly7IxPJKCPLxC9WjOWmDDf3DqcdUHMahVYb1HYg47YHIYtGXi0JL4v7A/ytU
XeoFPGGBo71+tSgshP9zffKAJABemO3/aw5YLnLWZ/VRF0u6/NH+M2etdEmKImuK
Efl5aX0fMzVlhCG/teqYh0UERH0k1tp2bOeATV28hay3TbY4Ry7UFNL0yAsUfjOx
gEdY13vzpy64oD/IcntuodbHJRSDcQVjuibPVW48yC4BGSTKVf2nETC/PTrfiCdN
dW41mpecvZH8EnxxLajD+Rzea1/pImFEFDtZgBd4mx+6l+zRIlORu7uNJsyJbeqL
/ZwPiJkGFN8P4b6MHY7bP2DiFf2w8f46PRi7CFVr489WQowdyPG5AvkCZanJ/DpB
AV9ksD7r1m7iU2tKQgy7+dAhppxeQu4yH7aPmGQozL6PB8Oz8KIDkaqctkD5EYIH
y7f5FMUlXe/OKSlvOZ3uQT5LBfne93KMGZ8caZEHo7ChsCNr/gQ6NN3x6Uzmc+2N
0anV59Tj1SO5PQTV24NmuSqjC20U/qkDJl5tU3wGnUrrJZSqZ3T9fMMdy9Yfgu/e
tslehnztoZaKbzweCLutFn1MTAqg4a2/EO5ZIwLHr3PaRLrzjqj6KJ37WIHN3f60
LSdUP5wgzmE3Hfzj5Nz9V6cm72ZnB/+GhA6ISnnUbk0LMRsKedeiq7A1yO9kNO5P
hC9Gbv+ZNE60OcJI3es3rNcsARTUOf8KViZRzGyb0XYQsbSbPT6wopuRuZHL289x
9izQ/qPIseHjR2sD59ZK1iQprT5EoP1/gCuCQcmFSm4caZJvz1CLhdLngUlHF+eV
sycS5HNRprHGmcLe2YXdki5Jq0nTpEzEQTYKh3HyGDJxKA/IyZcOVXH/Bo245hUX
37u2OTbKc+MiMzqbECG0dyk3VuRWUqqu+nGF3WH6NQiMsPc0XSPjgqgv0I6PY+fo
iX41PnAgKSdXD3SiRLwifuByvfc5q9Kaw1foiD2Y+uiRhZvrWUXpYPeOPs+0L8c+
urb3eD3KF6uGzD/MgKsGbpba7huTf41ZPoXS080RS1PZt3l8UAcNCc3561zPmcsh
cbmJkCMpng5D/xuUB9v8XUZ9wS/TtPAIun3HVod8I23D67jGXChdstA9y6ksQaFq
4J7TyYLzdW+/kqC4fWpQW9JVc5BwK8NYQWa+yHEn7MqJAWpq8nFAsLl+llLW+VAp
WVWypIjvYnlrtvsqNwVlPRznZRsm6H/jdrNKHxr3aSWdOHxOa/RaSB15AeP3CNxr
cgluNHRnM6nUF4t4o2469YFrfAd0lwR6l7ZicTfX7NHt6tHx//VKYRQ0B97kifX1
quUatSr0fsUHgQSZpRxTSZqbqaSA1x+OBsNTDgPzsW0kU27cBZUSfplrEWeB0mIx
JCIuzuNqA7LnuhDq/Q84y5gEihJ1LlSTfDpjwG/5F8hRnCZ8IZm9jBS6qgDhzIDE
tC5totrDilbylZYeEghNX1Xi7w7s+cHKs+EK9A942eYG1znRrggu8mjhohMxEtkM
j7Ix0OQSxvGjXyvtpJTZ1bYpa31zZ5dBHBpdvTptuUhUH3hhgUaz6m/vN7jP7GuE
ZuLZ1Co88Zxr+sFl23dveluTCoM0X2IstAXIsjrlSrZWVMfRFpySLqHLuYTh0AG9
vV8Eg4QWzqwa5fxjC/v+W1o8lXfKua1BNEIQY2ILjPltyH2VwLWWpk4PpsqRO1Ag
/Av7ZRI4lJepq+neMEyQxRlSmjjjn46HzgNn9ZvDsvPVB+QsEvwyP0g3SL828dXm
T9rlcQ2nuj4Awin5FPzNhtmm/MApRPYr3pcz1zxxw+vxjH/B+NzIMQ8iFR0L6R6s
mTbfnWatQLipHXV8zdEXKbWxbigzcSXq5+kctA8XpmsgrQCm3cR9oSZjaXEjZCZS
D/bXI8DdyFZUylKnhnxR09lS2UctWQJDH//puwzDS0ofeeK50pi7FN1q3WRaEONC
9ooWDm2lxZNv+Ax+SBHi+C+tTnzx+IrJ6CVmQjqyC8JJ5KB5N7mXFRXRCUaxTDSb
9VqojqxuoJ0Tqk2QnnHXlrHIbosGqCic8He3cKWbbd40JGtp2KL/E8Mssqsz1XQD
rIjmFZUg0NgAmIWOYrvKOzumE+pdvKzAXZ0HUIMWCfx1EAH2OS0HnYRgl5r+L/xB
QfpXeHHPz7yIAxnspqfmTrYAhj6VGn+b22SjnG+9ZPwbjaF13TiYrUWGtfZ/wUm0
DnGWNpwJYE4lEWgaU6CALlcl2cq/Kd5/AX076n+FrDh17ulFvyWUwBLCNs9JMloS
9G/O0zqsLa5/abCrOIzdKOiDn4QlrHP4IA6e2cZSXz7M+DAKkKZSnfl1I2ud3QHH
En4u+sus346o+kG8V8WpVgcvqAj8NC3TNSzefTwbnDOYTI2ke2fV+dwPjlefpl6Q
L0z4zWkdVpCoKnGgPOp1YLeKMF/wrYoaN42umxen2U5iMtHMnezIoGU8weqxRmYu
Pume9g5AprZUHJAta5Q8vych8NqQ55QKcOflV7d65v6c1vY6p2VgDxrxL7ut671s
QKm2IURpMB1P0wA1yf5whWcQ+Al5P02aKFoo8bQjr4bWijgyYXO934CHRbnY75Nf
YY2u6Y1GRLcaM0DEAqmyyogECE8Dj2cqDJ5WbnQR0bRPnTxEKQm7mTRnKc3JdKa/
SHEl4kknfEMX6tjqUicBO8hqSlh0gZvAXRVS5HoZiuZDqJotzJMyD1GzVYUNQZ8p
aOkbJyVUIVE3GvcqV1O+GuoYD8wqVgMxN6blhOIzWYj6sTjm3Qf3YSjUHuGeT3ag
iesNwQ8vp7MGaKMaeCGNaQJvQEekPqQS0DS+ZuedzbyOAzyGVUfsbCIEjYGdsBhD
wZzZW4/8mq18yzemN9nayx3OHInFyqfHzwKvZ+cj/CZdinWNChgPDVsZZLqKUegU
IxXH0IqPbhx/EJ7nSbjfHBf0PVlVcDNsSZQ8lVikfW0FPnfvkDs6yGV/CdXlgsjH
W5tF+DPd2hj9uiI72lBDT6aYOt69C2h8stOSxMjAPFNM/ujIWj3Yj5fs5w4lzmFk
1OqEYJMNjEtrMPrgx0z4/YUQe1GA7cf2ZZnWvdryTdkfGIQCO3Tqujq35PosaDVr
PHKiFW1GZCXyhAJQiO6JEM7Qt22sAmgiPFDU0P9Ve74b4dho9Cinl4fG06sggwls
LwH9mpZSl47nDvO34tdwTMzXt1WHdOlxndkKOk1ViakONi2eQTz2NH/RBQmbVW9r
ahGRepBmw67mZ0ZEqh2gYQ59YdLIEGLOuhS1cXfmttpKobAbRV3ahL5TIFqJskjn
DYWJJ88ronsHMMWDZ3DFnjW9HE0AeFqn809tPhP8DCyInNZAxunfKUcJiFTpoakE
xdSZuD+t3/dnbJVJZaJAfQa4BaRo5lxTXk3UzzEBmd2YUGFCdLhwniXyeGeJET1M
x68/DXJcCzMGYbGBT3uHaMKIRB/WA8gd7mEPX+ix+MA7EpBx5o8PDHJ0/lIyUFJx
XBYOU5VcoauqlPFRuTX7R7VDX1Zl+whDRaBAuBSku+w4VDs6XJnNTh5+3uIcYp3D
KM28QFrFx1jE8HA5Vz0FB66D/sefqPg1xP5ID2r8f9K3j2etkSXbTc2nRGmZYMXH
VuqUSW9hpf3YQ2L95JJGzTCB0QZ/XciyU98fr1YzzD1NnssBWqXsWPxQLHsu4MGg
Vzkyoz9F2apc7X/jozvYs3eiZWea1M4Gt/q9z0tzgbrXA9UKzua3aZpCOmZiI9kn
o2PqxW7yrBpZk+AJ6CVCpocbMteUb3ZnrmD7YMat+hMRuW4v46jdSEL38xXLfkw7
CMpOkvvxPXmzFgGQXXIeV9PpDEdrZyMl9JCRm/EGgkOybU8y6M55FXvuYjFKNJqk
rIX9Sju9oM/g4Jv9R0vgkP+a9GKxVo1+r281I7/6bOL1CyZr9cyPclYi9+xcvTv4
Wmbmvp+xqdml0aKfhc29n1gYmyyw7ivujgy3yBadTtad92GL3ycY1jVmZdvCtHiL
9O1v0YDysKqadfayzuSN6a/3c3H/iN6O2o9VbOZJlmBZJz+isO1LnLl2K2CGSZ+o
WOvC/VAopcJk4l+5E6sKT5r9zSe5cGI6UK/dfKbNOs4hPFCSA2TBwjQhRUZvY5Hs
IZ6AtM0wxbcxOwKyvvUycoklPU72hGznUw+2elMluBwMOOss9XunKN3KZGrdDn4n
6JP0fPiiv7foqtbKUUYRtnyEsANoeawSZI4St3vR1AVWmNN+uRW+QJvx+ZHwpeVV
cbuGf8tJqZL7STUv9exjbyyFs0WSGQ3oDx8qLKxjeurFZBkhdlTc0ZHb7ouIhPZ/
Ipbm0roVQczEDNvYdiWm5VordBf27Wp3AArwtnGQcg/nqY+PV1hSDGdRdedXaN5M
veXpiiaulqzniW/YA4T3DIi3UaGdlWyPixDD5lJR5N327DpM+F8cxKkLOeAT0jIy
CZr7DRikZASm8JqMxEO6qFUzGjQzu6qaBj1dIuadwhpD8HcVqyrfv61fDYktCe/W
vG/SBeGPeffnH3xxuhcbwA93cR/N9+FbvyxYqvqZuY1ypHFDBmlqO8MLloWzgZzB
KsjJP/s5MOhuxAiDKMV6fQuBUIOnRAS7eBGqmymucctaYfjVKgHhAzQzNXUz7v/O
cs82951efFIXo+Q2JFDlN2dUDzjBDJ4zVCX+o/aRrGpnn7TcncNU25/qM8Nm35e4
bbAM7sf+hKN+pWRzzuHb9VSYJhiBlifuzQoMH+eX7vF6q9bQTpxImKVA8ocHx3JS
ynCyegTVEzTBtBy7SE0Ob9cnKf/L6XcIjNN5CVpgIvtPLf6I/ZrTVIQjyzXz71XD
dlFnaUB75Ke4C0mg0FQD7g8VB6UWg0K4dlWyYTyVGxNWMfCeQLyEVOH9IiAqQMea
gJenxdG+zkrhI4tKL0S2EUrh961Ptoae2rT9HLAoWQqP/+cyaVwn4321gebDC9uy
FZv63hxulqlXZDkgSoIqutfGM6OgFpqd6MQI1LTXL5T6we+IXa91OZI0htwxYm7X
n9XMbmrRuNiIG1w+BgiESdtniQhsGVc2/r54UGZi7vaptK8fZyYeV7GcNj96tjC6
FpQqO0hPh5BN3RZfoRb/LEbs5V/J5Soe3mBzK+umwpe+mpFLJTQnJYxYmife3bh0
h0D10A47tnZjCFHPWpKDztdn0slm5a3zE5t2Zxuxj2Y36vEEh6GuMglRfwkMjf6j
eflWNsx+DU8UMd0R3ohWCHdi9wkHqrVreDzXy8791Gv0pxPoqFz2thbAB79j6ZCi
9A2wlgEw/dsHqMWZgd7wl2DGWtDlEnXZI53y/tY1bbjK/P54apSflchg6uZjl4r6
DGqKVeQvQ2ulCeA4mAZyAYFJjuBKyh4aUQDVK8sRgTM5MOs1PL9iBH2fu3qy3FZU
l2Gtyxwn6loA1Vmf2Yj91mwN/TO3XOcUyZf7JmlfOl8hfJqhP3j/q1cDvpPXFtGW
2wB9/O/kUQOD0JF0p2aOSgD4lVEYXaRg08yjhLSzBLIemByoJm8elG0JeCc9zGQZ
C/bo1UQph63a/G2yyfOPPHoAsHuhcZlypyRxzaS3OITiF+ZPPy2I2cAPTM/P3Tln
tckDglktUVf5oo6wu163nV8I8WJTGxrS0iaSUAaWi2FNFBpQ6jR4nCfr9F9DBir6
m5blNsh/YX9E4uhZvVeWmJeh8L/1F6gsUKTAvaM1DO2G9Csds/bPI1h+wlhszqdY
qNLdSi9MCNkflFPqS8sCs3j8+iQhSia4BTDrSjWV/kAN2slIp0YHiBgDzVieZWNz
J+aVXsqoCOa1NsadZYKqc0wlMoBRPzZhFQ4bKnbYFfyhSustrr5nlZG1Slnu7Onh
apUUkIjOk4r21JRnj2Z4Gch9Grj8f76Zvo6KaAdOiz000ew84JLaANStmEQZWNRR
U6lBt/s7vnzAGVuqFnAOF8xaZulb/V/drxTJ01HDY+FTfjGMLFg1lopo73K98Lay
UMExCNXgtIHGG/5iA1E1L/mZqu6hSRNo7TPIaf1z+bLLDhBZ+hG5t3g4ypWPECmd
P5a2iLyMS9pu5yjNKFw9gcgzFZh8GjIIBvbvMThkmoMTq3pfqW3lSNWHkJ9sCMZF
cGBXZQtYOec+BMrtO431Ioe9qXGJ+AgxQERjb8SaCARHLHo2/Nf8XHP28WWnZyC7
f+8NqBMNIqNrftpdmQTOFAP/vQHr7DAUa8BBWMxShUv26IC8aPcZKsL7001frjOZ
YgNTlmkY3AypGZmCJ6UYbcgUKd5fBtad1QMp+NSASKCZ6RCX9wvDMkTb3+8uOhjX
7cWhmh00aQ2B6vyp+YEGRQTFWW+TjaVxvyRm6j1b9L/1higeFIkjnWzxxWfEJ6PT
/Zv31l0VguQOBTbKGC+V/wfMELFz0yH9Twgd6O49kHM4ZOmMZa5RAJpYj3uP0tXG
Sy2Pz5YEzQQpHG/EtVdWysclhEBRe1M/slnXaRpnkvbEHHkiuqm203rKjSUdpejL
xxhls7zAmRe03M7vecCWyhkNpJmkplcdVez7Rum7PxXo84CA1CeZw+irC2/S077c
KCFQiQR4WO4wuxa7Pltn3F5YfOzCPiIf0fnVkt6Bj+KJD5699Xl5lYwXwOl4tGu5
5/Utn4u+y74BpdJRIxh2wSEsLk63bQ4znmM/tluxIRgbFeMxGQjxtCTMndPoQ6yS
WY8GghBj34lmmq89Alzx48QzFpYOgYnsI80lUcUYddtOSLgSP1h2dKPcMcpF8SOB
53i3pQ0kMkmdXi2sGWlA8avJgwD7cat5kfVQJLeCRUzMXaQ9BueZBcQKT0lpmvyc
043VfkLunmrEahqdszWdAN4+dZXaRMxJn0Qtn6ILXrN8ya9Vvqsd7hxt6Zhl36we
fx16UO652lBuvNFQX9v8V4Nxji6+H0YjUZCJPfEp/plMGA+mCj1JdMZ3FANPDhpv
vCFxkPRYsrS6SzvUyjf7oCMdM6XjXX4zkK5d9rRcL0qQTsSivDR8XVdBQMImnzhq
GqhaS3vcJYMwKEo9RqgBEHUdVktmueOyABK+m3RtV1llvEJP+SyXeVIVUo5peqHt
mjr394BmDOanflB1ZB7qKGIZy1oWb/y80sF0kWOfZL7kqtucgNObavtvI3cAoFh1
cVryRZaczukzR8EUhlZ0xOVcSNuVlGBL8Bx2oevI1y5KL55PbQRPJKA1lxAYuGkr
/2X3QX2M7JhtPk4jgm5ifSTfeAv2e1OkteCby1BA+Rq+Szd0T1q2WFhRh/NKWPCA
N5KFtmcCrpzeRRQdFwvf0SRQLB3PEWlew4lrY5ROrwYj17xKPRQ4simlXfQR5Qoj
M16FgS2TWAjnCLfCzuYS9yy+Hzz4dMnFpfQTfd5TZF14vOkdxxxxpjBuz4knHJvb
izVotdLhtKgSgji0bLXK5wbN+gsDeYgt3zJYPxMeQ166gitkl6Iejt1hK7hl8tmd
iY8U/GtdWgHHlL4ke4TOZQvWP3HAHjbZVNmCbNffeEByb4Jw5AVta16ygMWLDN7G
9UK+BBvpPGTxhziIX2QIRtwEbvbniKM3VJK+YdRU29i5u4H7ckbBgRImtG1DBbl9
JX01yu6qF90bXNnyftGvNysgddEGgtpwjWTsk0WB9Z34jLLI0SyOcNVttRkRAmsJ
eEot5DdMYzFMYDwci8LkC/VcvR4F6FJEkVQ4sOGOzMwSkBjPORhdxsqWYbAUhQnP
luFvwT3vPRiawom1ElsmLtsiowFLrlnGeXarDq0FrRGulY/l4u9QNyYWAxalG5Iy
gl95wxFJPSNp+q4UMK4J4YhHWBboZ63LKuvQKpk0NSOlPaJXdWP4E1PcDDs5wxZ/
S0rt4FEZUE/qERsUh3fVWa8bYTPFEzGB2Yn1aM/UmcjaCgS0vxWi10K8l9aa3nVs
FrLgguzuSIbkQHYZfZZbknibEpPihKF2rhP5SfvITvaQb4swadFZaRMCc5gg+fwA
u2w5Uxvl2+KYCC1Ti212BzjvdVgEbIiBRuZiNjFl22I1ZdHL946qHdwzPLly3fIj
1noxhdjh+Tas/N1gd1Rrirg69+Xbki3/Y2TdognCUO4xnoZSMvpyGsMb94WjYUvr
fJ5/qTjnQKFEJQ0lNI0N+WXVAc56KQ2b6NKyqwsZFjCCZzmIJ4sD4B1ZmYDqXMvd
RRjgtnYIJokkYH2nCVs5mpqlyIpZoH4FrObYK1EbVX//WWUy4n2L7guCLTcfl0UB
UsZlct8N2j8nG0vmsG/WeA0SGBF2UfJFAxXoSUv695ThF61KzGOpYhcq505qBomg
yYGBihgB4Q0yDMffm5tLPeJ5Cw1LuQTyF6sqxE00AoFhnzc3iv4WKycG29JBrs9m
nsDb3O1e/zjYrapMXwIYDiFjYNt6vfPh8ySJMZ1ZWu5R1WXpGom0RhjQlaluHE9f
ge7vhUl5TIMmNOgs3ANEmxiy3/jFRzWd14RmSatkksHjA9RCJ+QrMnt1oA973m7T
oVvNGbUSfoMJc+JmGMwlpQLtF45uri1IeuYsxAqy2hWz6wo1tn4iyXike+4hUFsM
+yDDEG/TQWlHlvJ8ByzOCdaGCazU1/SqAg1QK9D1t4wA3dtapx3ofXCkNReBquNA
XOPKKdx7mEC2W+njCLcsm2KB/C/9RJBiIfpDD9+81CQ=
`protect end_protected
