`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
A1CCbce2VJiqwuIJnx42WlFi6j7mfo5MiqBNC1CmMvAaLdECzPrP8V1uWRYpS/It
4tas/qeOTb/mpH6z3OpU5OD7/XvVhZn6KtgeXYsG58zTHBkfCa0vqb//bzl/19yj
QhgkwHcptT3RVuZfMtFLqgdL9QTMzRRseVqspr5huoipCDX8oRdmj3XOL4MknVIK
KI63x2VpzVTUlJRDfzGeN8UvbObHyGSYx4dvmSUmsC619n5dp3UP9MvEvcnDGZsK
uLaYR/UBd1u7zLX0QwcogoXe+8VLlyfDlv+FF+ggiSmGRnDACeN2nCMc9gPeQ6wb
KT4RSPERqFK9WubsPFCZ+Q==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
UyE0nFDrlJGHQXmwcgAdXcpNa5YFv9AbHauQqp3VXtFeFTvFZ5T3m4KpXrnaG+Vs
wFU3BxC3+JnwZlADZmDtpaFUMH4ouvST61Zt3n9xmHltiZA3vpkEIT+2Or5cZfoQ
mn81puhV4+VVYA/1jr7LgzvqOAJgRkdMV7lbfred9lI=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`protect data_block
VJpYeZDC2vU9JL+eSTG/lWbwyiC075s4V+p3bYWTnG45Yt1ha9FpFZIvT5BRbmmg
JnJ+7/y+H9/EOPkD+L/fX8kMXxkdpXDDfgD6RwOUvx+RBiqNFvIjpeNj46vCwdlC
4BFdaD4zJX/frBeIIAGf3Dl9B93Y98mNDvmiL6BMFpOgnOwebyZOtQ810wemtboO
89IAqfri8uE3i9ACsvTYpKdpRgZX6+jrPsOxIIurzxD8g8eAal20Sik59bwagL7a
yqZ3G+UxcpcAfX/yvNGEthCCgrAPbIH7AlSFAJnFOW8Rv5m47qKSt+9qzl7UDNvM
D1YU+ZebUJ4xsGeMUur1H2FHBZ5csfJnChohq8LNDIlGOYjjChWRGY525c3kNGbX
Wqi1ixYWAvBRsW6OTsiwapcGRrzmJQAYniBHjJn+qi/NX5rxVh51d69sCxdf5jpc
Mlxoy8c/zhDfDL5K6disOdBB2bvEb6ONGYWQk0A1gEzj87kNcvxqPb9iBupFTLOj
QiDq2l0uHReWGLbdGGG7Rl3mNe5pkd1OB+DCOYMoOpexjJB3ba3iXYdm0N0pfBuA
nJFw7FN85c6l89cE27tYWYVvdDu8JjSbikQfpzP+IxqWRVBZ2crVunI0qI0JsR8l
EgPjCzSHeiPQG8wDD2rMD0YASr/Gu726pONbQu/EV8JEJfjjzk+uC5PFInjr5c3E
yseDk3tZPnBFURyvbdUIsyGK/fmhqjuVdhsgBMjIlGHHYJDnh5p35zFEszN2C4CA
o6rSbLHNOoQilrgPp4a1k/9aC1AHpN3p2sgsRkMf07gn9rLqwOgsJxRlkTRY1dKb
yKI8J86UOrZz73gPKVIQ7DuZwlFsJorQQhCbUtvn5+/Szl9036ZhyJDahACjh2Fo
HKzrelt+SAcIv/cGQmL7umH8x/ws3p+S+D/vODYhRN2ISwvW+7cp6NZqjEvAX/ds
Ce4OTqT9FZzCv+D4ts/jadrA68Mb5F1vLsJt0z2GV7aAWCStfqwksCGS6wJFgGRr
TSXgT++pwC3ju87ixz1XTSeeWfzWXLpoZoT1ajUhkIv5xCjwhdig1+JDUQ2Mmu+w
YcJreGv+ns0fr+TMB46ErgmlW65VIW0iM0l1yoNmDjjk7POxNCvzMF1vSk3lI8T4
yvnayyOcDlNUthEo4K18T+i9llnkHPfrNk8tO7MQTG/OkjDkteS8jVNrTeuEcz+X
UVpp9Wd8tQBBePJHJkXE2qwBk3uF3LLCoV+CGHI/OIOKDkVkLYSGpgbDJNr7PLXR
vQkt73u4lHhnITi62uu8782tHGcGChUtFPy/0y9Se5nJShUQjKU0UjheiNTfo6Au
6sPOfk57blnsG4K0Fdfe2ozJ+2D4hK8SOD6ed5kp6GWdJ6gUBZeGRrlvm6jgeU4m
BFJ5l+DGKCCWXtaW6tZjtXKqLytmY7XQS3hID9zs+Iqzt8ozemp2gfcajn/Yg4Tv
xZIQTjxwMDCQoJBEVeZKn6koLW9i0sRWiWkpw7b6usuVfBo62OzNiDDGNAfvGV0n
vjKzFul0xxjOTrShMuwOcBQ6lLSm5qEdCVBT21Dr22JD5s/mADvE0+IgRFD6OYyu
15HmF5FV3rBuBHoIUDL9QVdfYP10tG6cUulXnz5nMkGB0sZPY/7YVMqK+WjDO36q
NWH6TZTGggn5lLjgF2G9R1j61TVn5fmODq0sE50MzrOqZXr6rPejTP/p6VuCLCY8
OZsSMYiK6VwOzcLx4DRcWiZ3DVj/hF2e5KgfJNlxBeskrA45V0k6uo3zGJF4fPsk
yS3xxmGzxKyxnvo2jo0MqaYed2ib1chrG6yYBLL5VWMz7y7GVPL7ssThHFNvRMGK
AqjUD+TZdmuGGPqBAco/f/rcSRa1zclW7Yi46yAl2ZqVR2KhTZiucfPhBhr4thUY
Kkq2rUaoqPOxf37DIzqAiqilCrbQaSDynVjr80TX6yn3KFqTcY2K6LevrDgVXeSI
+Th+XcYRyKBv/fm9kXSNjtiBPAVrxq68580/zXqraiQtRL5DMA+oCkqJRA0qGJHy
l5rwxUS5eCMzBqu/We3Bfylv7c0oODzdQ/YFxSuEhWIlYL9BGhOxjQnoDT4Ry3w7
mqVCkElWVeMFD9YxU/i0YOfFuqoyYXmeLhOyCCdicuNY2TY0ZlXGUNkInBag99DX
8JkHJkN7SnZRhSJQOkH3/Ptzh7PQaEoDUUxoLP1KMA0C9i5hyhvMhiC16+Alspif
vHSsnAicnoL7TfZ1+0EzDWB5/n10UwG9yL3RcGocPgzC0VLYaSOxXltP5oohjTCd
/iFA6gVJ92tSp5NEUixjgz4H6xnssVKaOwLO2s7+8cveJGdJ43XezQALIjnXf4gd
R7ZzOLG5Mn5HYllReH/Xh43w0Buo1u5+W5Rd7gNtul8Cd6+doHkPrdwCEfzxQnyJ
FT5N87Wgd4Dz3KXLfCConmWaH4icOviU7uP9GfYhSW1hV4GAlIik8RmOu3b050a+
v1HrnFpcgrl9vRxc10/C9Uafwq5lZw3rlJmxhwAlzSFcwfWMbBA5/RQgf1xHSpsb
cx+ayicyh/U5NXq/QMaSYerVR2GxVMFX4d+KgcK6+73fI8Ds9JhHWLi1mxjY/scU
dioUzc5rzb04TqekGoB1+mkxKvQ+X4329TT18BcwvuYHAdXvc69hgKg5F3prZ7HO
1OQLj3qrP+5IeFyD1RAxx12Qni9N6Q6YR8oouVacxzCyzz4DkU6Ojcj1uSki1wXN
vMGCTpMRZimnB9x2IF6+1QwNXdzA/WidBmAdJROpUksjHbaWpL0Y8i9TGXnGB4pl
U5+r6XbBuaar5eScIr486hQgpaDIfZ1qVKt9hEXoQARUf7CA5VjSxOItV1r7bbgo
z4BH+cXI5gc//ZkGMkBzu4JcfM1k7miKn3Sk82QrRFZASt067YYYL2pJ43wsfrYR
sPOBBESDmITKWjmGz9+mexnIGJM+ECR59Q6M9ZvgWerYQ3+QLK0MRITceR/3/jLK
tarYqSf1yIMVePpx5B6oGN0FZoOxrlwTLZxsP4oewOSpsmK17PodjewB7OLvClVX
6zUiFVN2OcFR+UkGSRLvsXg6VSj9p0OqbmV8TQBVg0uxygIHQZDWplLNZKgrwWqj
EwUP4aYhL1XDmMCtKDBNOAlYiw00xpa+6hSw2ZOcrHtn7PyBUcM6tXBy0uO/3i+5
70M73tS33ozCWyOnZanFU28vAsOCCeTOeMK1U+jbmCjzhZvhlQTAuF+v4yfm1xsC
pF6uLZXCjoEjidKvF8Ju33GzGoUNg1FzQTHFp2iwW0dqrY3w3yggPM5mbfYmGUSm
3XEdU/fDO6V+ap4fdSMYv8MjPY5tyNWrNu8Jy70tm1O2HpXZRuANKqMJ6lAyzNqV
a4OJmPac9s9WVz1hviNDAubKGMyNd63UhXIxPVLt3KZIuQ1fzpCPEmmtVWCULuT1
B0ICWPVeUmcFscK0l9ZhCqzww3ugusO4zJsC23deRRbPD50L0PCxyNhxlHEVEepv
1dc5pRBBFrXrlY5BEfhfpotqqITRhnSlWLrdTceQfLfIsq2RrgIxGfPaTD8tm2de
H/FOFUJwbDWbL9R3ADf6HUT4qvTLTAlbR3XYIknlRXf8Fcvp8x014KbHx2KZPCd5
OQVQiZfD/8cszuDUuE8LJZLg0JUnDmyFCmZ6gmqpoZwnUrqzSYykEqXAg4njyLha
5GnqyHvkTLsdCL72H4sDOlx1PTL/kG/T0l7kgRztYUhW4g6Wb3a/lwj8QKVtYZxL
7j/3/HVLvRLf+jzRegs6dGkcL1JFJueclEqR596+sLeFoJTEw2mkIhPWLdidSd3O
xlgMKcHznPcNE3FiAKzPae+/5z8akU44Aa0Mh3hImdr066HtvO7H3R+WrOyepxKO
xoDX99azcQB0i5TyiIwZ2Xiv2dB7UwyK2R3k/4UaZW6lI4sIFlEEfKkrR4Yyhjdg
L7uyNRj/nYAW/wS6nkqqKgBbMk/TKjgkBUnND7PHqapaeqIQNQNQnoTIjEzpwQYR
LzTHSmB69P3DEG7yE4KVOgly0yXAgGp2TwS2588oeB+xieQ+YBHQd/DR/Y5WFUud
nixCwenZ2qx93jVot4NXy1FZWqjFkCGLmxNxOzDkeV2swDx3QWwBKi4y75USXPPL
VM3dnifqH60RA3Juxo6daSnR7o67yzmR1cYOEB+tUSFlgtdqrKUQUEVmt6m85cN4
YKcEMRDiAtXcpMU+weFXOvIjh/Gb+lM1h3GlJMqm9F62NJnzz2Uues9GV92E39mQ
Z2VipRee2oSoZ6jrYwUhDWUUARQujFcOGAtUfOIIn/NeA9C2pBLTwOFYQKn7Ject
BOo1AgMTOY2WQ1AlmhafL3bNSzeGSOiHe5Miy+ygCUM8/HSTr47HM53EodbMhGaF
DhZyMC1NbpvPrboc9P37l7sopg/4DEEFwU1cDqinVwktU23FeI3apn+Gb8t6O61+
iUfQU+ShogTQkph6FQorfEFqnDmXl95nnI8x/usLsvOk0I0VS6YHNRrPC4DaHyky
mH9hgK95MjOyRY7MdmcIiMdIRdbH+Ce0izPJVbD/5llvykhPYdGvEffuI3q1Tl48
nap5D02pq1FJlqHTvu6eKDuPyMz5SLDRbUxV+RoRXIVmNsFd+cJS/x2MmV9THm9L
IbfmB3+Ws9QufShYzgbYM8dUOLB1MJQ9mcqoGfD+EzeZwAlKCHI7mS2yn33MOTaU
ovSzTkwWpr/d+3UQkdvk6QqIwr22X4zkczNa5rJdUJjzjXExLXPHkkSTpen++5bC
6J27C+kkLDO4+tATLEtlYEHcD9BymtzJJwgRM0jbyDWObvvWA6CAvSf2sX/g+U/y
K50JZX889sx6vWLoF3s09j/mw5HBABztaWCkUwEa67/NyabP/bgwyrhR9PlEYCYA
60IeFnaStCANEDjp19tBTTsrbL9fy5y98XlRcXhhYuen74YSvX7dka3WV7MnY42V
lMHEk2IjoyRqzFBpljAw9eKyOUV5Q2ReEnDj1IV1QNSBUrUBrAqNs/V/PocAe6qx
s55XKAQ2IQeTUaNpY1LMi9yzJ/x5NgfwdpVZjT/V6Qfd//KeVvHlMS0U20PwfomH
m9O1+tMfmgTkUh92uFMvIF797A++16GxLQgRM/VUVbu+Z/uK7SpABQUp3Q2Sw0+v
rp3mEaHm90pdL/OBa4wTU3ZuENNSqURKT9Z50ATn7+MOYJJzoOyhOg45T7w3x8HA
PbdxcRcLkFHdtU9UmbbALJR7IqtOn9rheXmcBzAbg+COvAYrIzWGe8xwzf9H/mRb
1GqBXMySh6NNv2kFOYTmOCZJqsaj469QTaeqvB+xqJWoSuIw5uDAyljOPReOX9cT
In8N6HTob5coVpVRfYGYqw8MHWaGTmYkjNF5NOdiE5Y0W51ZRn7SMK1cXYGPoThK
zvGkPfFMVvfPg5nwtL+ILh4c/4ZcDPFERrj6mqMNh9PTeiAEuAtMH0MAjYcKVhMj
S39iQcZexBGn7u5kDkmpo1nRir1u/wDOdn6k8vL/LTct3IdwcEFU9X9OBnNJSO21
us2S1p4RPY95bpHOAsDaPtLvCRgWuIWZx1MgeuIitlOoPipIEqD0YmZgNn2n5Qbs
WNXnlk/MUrMFuA1HCIYoi0fv2EUYGeRvpuDnP6dwhcqtH3rmaX31DNx27b6BfrXJ
Edf1Jd+xWAu2ubqVTGnVL9IFpFzqgN3jLX1YsURYozcwz71Sq8al4sI3xPxFyGPE
tYaBDFhMqnxQsEJLuaYJ11zBwUUgoTNYysnZd/JxIsSM/odvVw7zIrJbZmD5wWSt
Rb+8FwXYYnRJ6OJqyZMHqiZ9z6HZnuDs1sYgQDaGzZTVqTDXHzBVw2ewvMGnNXSm
fiIwL8q0WkKuf4J/PuHOhPuoJXxFOp4f/HDMOKP9foxLJAI0yPvZOOllDMZ0+XWJ
hiTQgZRfXwsQPpja1TD4uhZmNQv6nClEk+YhBWLCXgqYH2AhEMKPrlXXYKqefyhz
yIqb8VvXfMX50n84qg/q8gJVoEIrMJ0Y+4SM544PI+MXAPd+aVv2an3goDR9LjVW
6waWVYGyRslsWnXg+L72dyd5raS261HlqYXhtVZ2U5YQub8zXHZHjKH3CYdAJ5pl
IuUk2OLy+C9TipI8fH3r3nR2fvQrewhRVLS6XPxXoU2ayBkXgLVQKxZAYkv7HzNC
3RX4HAQtSk3Ev8+cWf1xyYWEXTzVVI4/S5a4YWOlXB30xvPOYxwk84S4+603m+Pf
A/XbThOn/CLLgm2hj85uN/0X4sCUBCTD5i4ztnRIwSqnJJB4lqMw2QWHwXzu4niH
nQ3vfEX3vwF92SeNoqvHoEZoEUVy1UDj2UwKrnOgumR+Gchx3N6iCPH4Tunpt7+T
1V+Y8g6XIduSQANBiERoNGSEfKFDlNF/0mxMUwNLt4+MwZyEpJwMItdKoEVdUEC6
03TLyNXHu8YktmsxD3q6m1u5BBCBLpBCqnxGXdXoU3wUwk1Bnms1tcQs92yfoJVP
nAaUOJPOmral3XPJnkC2fA4noEZEXQ/pFSLgq7YTkItLP+e0FbmfkBrA72r3Xmz/
S+ncYREeiI131TjitQszJlu306u1B5rdCcCz6DJhsJo9niBGYoasFX//czcu34vf
AZpOGavUVDMTOYE/ZtNOh3WRFifgCwsbvhYn+dTB7nPZGljsoNEE0R3NcOz607uf
gIBUNfLS+r59gxnsN+C7HCf3RHCPi4pUXP67NqOdlVKeQclApsTTtKNeLZWiryxA
Ef10fOBB4LhnOpk2zrELIdlb4gA1lDbtfL0tLfZhJRBC66qN4JO9Lt65PSaWozHM
+nH+hZWnlYmSLYVHInIro/7k0WEzWKVMMNvpU4HV94/YkHcy3h4nK6iJiLnYKh7y
qsaxvHq4CLlY/HjYY7wTOocCn8Qt/gPdvQQnPPPskXxioHqU75F4lbugvItdAXec
hs+0RpkjNvdhNIITtfcTwU0FoTOTjdkObKVZmyJvpCaSJ15k9e6JzlNVSrRhER6H
+PyGgfT7ETJL5w7vCYGGjwvC5CSfLZbkBnFJZ6pOXP46L12svZn5Uu/RxFwKeA9U
bnfqOiUnE9UoZb8s7afi88Jmne2UOKC4JyfQJLp7IsBTVHijiKC9NKNAkQyIcNab
4ooc9XtV+uwI2Wu9Uthfyy0om5mM4FYDfxXiVZYOLMTvfFwqn3y0CFG4Hm6GDsXn
8tBcvYLIetIl4xbPg5H/J0W0e5dOCKNA23vF2cjN+q9semShTptg+/Kh1HHA50Jm
N64Eo50M5bW7gLz1IEV+sFp2JePUVxpN5J3e3BYWh75L0OqpJNVyMOTB8Y9uajbr
iNxXhhhPRyTtYd3eKUFP9lFvB6+rXUsyDGjMxc6ZvD9mXM2VSAsLo0NoLrk4giBf
ponO+wTE+wXrf693o/uvxpvCxOkx48Bs3rzIbweLl4BTRbkvbwvjOIhW0L0bAHOa
baYi1u1Y+r9tNXbQrWQz35LoBFthfavM6pHF79A8TcgOPV5h1ajUtzoJftArtvxS
hEJPjxC1rxBZx0gKTJf9jSlkbkvIRvFyCwptVuWKPI2Zd4jp/4onulM/X846Y+dk
AUHt21bOjtqib8MdGvdTHbBtES5LDhI+08SDDNdJkAhBTG1UFdsAvQJrTku7m26j
VmRKrrIIoyMLYcAof2ThKNKl7USeMLaQ14hIVWrQhiL7ua71x6lUQ++PoSLJIilz
JGj81bdCiadXAB+9N36Q6fu8844UoxTjMGfw3dvFzdXkV8ACzBiNydJ7D69Ffr7C
XiVtbPe65Kpc5VBWltJV+lVQ1wUWNRIXVpI9Fp0k21TIZNv8JTatUjnC5BFqyXJO
hQVEsUfByMR+Dno5N7lne4PBVowgvWN/Guc4JnU0ShYYUmSxq7J38Jt9nGrRq1oq
tO8J3OsCLtPk4IGI7MuhsD1eetXHLaqdt4gY3l+m6DBbN8p5s1le0vtXwAfoDJEK
9my5rHZJ3DfrIlZevDJkHFIVI3tb0Bsr72Zjwi7t8V7qSlWqUHD72suwh0Yc0iVZ
ssfcmL0d7zshE0PRxlsvBoFNO10BejbvKVsbX37nvLHonAXOKTbfKY5PXEmy6esS
V4QS4mC7kNAvK8Q9EAWzttnUfg0oFvVg7EdNmQ0FIhc3GE9uP/fq24ldKARtoEQc
zizXNzTZy+yQgd86px/6VZ4FivU5F3f7880lCeiRcDmXvSJAdbkMS1N3lxfSK5FX
q0e6YfDGZ939iZpW+oZZg5FQWwRQhcrxiXTHKExy3O7J1VAQeZfvjucCe2z9C/yl
HzBAOlMGW6l17ToxEVCbBV51JOEyI2L70IG+EzkuYTbO3fxHNDAzF/uwpKh685Aw
jcvQsR0MS3PfAYkbDQlzooQP1sQpnGDqtCkdCMKwVYs/y8gksshdCt8K4SQKU138
M6kXeXjR9gRV4Hn+xBi3rVLUzIbu0QUtHX4u8iX7qj3YVRAcjt7oSp9on+bpXty2
oJnIUHkdgqglYxais+BO/uK5YJnaYuYL5PkoQn3Bu/GmnNmol+PWH6dxLjZD/M46
HN9Rbv49SbA0vYO6DB5EwbhF4xDxSLtzvfbpkDis00UUefsC19xnHawOULd2BA4L
pYw38kTs1HT1iT5DTDfNqkfOiEBxLL+QeVvUWHrJvJn09xCHJ/ZLZ+rwQ9YG9MfW
UdCr/uz8B8ST3gtrNzOLUWg2i1ZIa80Pcv8epE3KPpEW8E1Y2vUYxfWYdygBmgIB
79W6jTBTV42kT1d/L5V0OSmBV6esqsC3/832HIbNTKY+eIFB3tm7Ef36UdrDx33/
6RvWRPXyCDePYv1usx1sO9IHBb1omFSrA8oZbXl6VvwxCF01JkdLT6PuVFd8Wu4y
KQnvzcRNtKOgb7dLejNzZOT+QFnk0eYQ3vNaxXbHP3P/ku+rn4W7UlK/iDK8tRgk
4vnAQmk6+4KchVhmpD9xXQ/VwOlWpoL02ixf0lGR37y1khZM6OGLNaG+67r/uYsK
LSdRFWogNsf2Ft1ef1rOIzlZ8psvHV4AUYvz673uTArsNKPiDm4eiZi+HD/Wk4Dd
skFBOcQmKiikv2h3vV/c7P8iVkPq94WKCXqnqD0DkRIcm+XWsiOM0JEeQ8TEh6tr
/UPN+lBdaD10khaXKRs5dZwj0xLlPeEcDv0IbJpSWtYZT4sPmVCZAJ8laMG1p2X4
3n8jV4MfhtPJDHqoCj39MbeSQItAyA4FuHtaE7J1Q43goQ8jYIbL3a68l4FAJdW+
SYn3lQKM0hV52KbICu1CeOoNb4pbqjnKQcAcAYM3uwl/DvQVZF03ebeOwrX4OLHR
Vb+NlmnjPdLlNFjtb3ZitF3lEkDaaUb1EJSyQpYTpa3iNE19iD6YOKSqYuGXHvWt
NMBKtcvaNSfaz/JcNzAT2l9pVUraBcEbtM4d8ylPzOUsiSTFE2fClopZwRMsRN23
GtcHY3EoIwiLbEGwGDnB+vE++jl7RY8o9BWYzsL3qJIz9nXhkcrLuUY6H7hc+zEp
XyaakezwL5R+w184yst2fFtJMobZpWC96vNMo8/M8xB3Jmst60ktqnFK3PTI84Qp
wl33q2kd3e3DWwW4tFnVYrzTvrijvcZkIzNMgFFXXJYfHIep+n891PLdHtStrM2M
9mlHpsgjfYA3iIk+M+GJF8OCiQ0qsFYRrwzm3vy5mjQYrJlBPrhv8kheanzzgUer
9g+p6m5dWOEg1v3MhOz6tEQgOzwObpOhpf/VzFqUk+LB5dG+Ba983o8tK+QBxAa6
H3CHDZmOdBOO2efz3wqsEX6AeiKok46SH0o452oHSIUTo8jM3J0e1LlmIg6ngW+U
bZGsd1dcFAI1jNxqY+OTxuJSfKJpzkb5E8CMnsPPLLzHJKu9R3U03ZQwXFFxDrww
prPbut5p3xpwB6YcbAh36JrU26Xs/D7LthOaUjEwRy5WRjziVfQWH/qFg7b+HuCQ
oDHUjqxJhBzRyAhSegpZQhfYvN6uzGwwSJtvE/0i+vHnGpLQ0rQgDP1JzX/VMXyA
C279d7mcbzI/mEmj7xBSsOyFMiUZ5jUEn+EwqcDXNA3VYe1GErYHuoi4G1LuYISl
o+vaq0cU3sXcOg2Ui4VhhCtPv2ExOt29Sb08EZx+AURkbBkfZBXAB5rE8UpKwzHc
USflSTFeGF5VkEBBL6hRzoIPiJ3mgOgb1GfcUGrM5qMUPRvB3i8XPk6BPo+lvvow
Hr5LDnAqIOjZtPR2XCsdBSwuCyG5e08cB1OhZZrryOszgjS3+amri+/GLMfVveBM
Rscofb72p3WfoKKJUax+1hyF0v6C9Z9ECZwlapxwhTrbUriQDI+Pjpv3WUtYTM7z
JDlh80n3tUA0zWU9wrJwzwxRlpzIWHhbQm0RBTwuX0pWq+CMYB4axPd8ccTqdHDA
3L9LE+1X6/m4iV81OST82KS1smU2FAvsGGjopj+TlRqgy7ZWnWlU/qOYug6YzbCU
7pwayvL9sCBLN53uLnvYGmAG5Ueo6JIh2gK7eapA2yTnyNC42iCD4riffczj2+08
EiB9ZrAEGFRz8/1j+AgotaHuTO5nEOhJXNNeTipESSbQxxQgRhshx6jQGCHC3TII
/5l6DSadNCvVAvbqDnVpx0EsL8TbyJ7MAopy/8pnXZTe77/OJ33EaZ36+T1x/d8p
`protect end_protected
