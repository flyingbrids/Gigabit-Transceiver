`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
T26xeWwnBZiSfhp1qeV/JPUQG+yAVk6K6Y7bTSr8Pl4j9A/DdkREVFOZx2r/Int9
pOvAjmXEmxhEEoLXp3MedDt44WvSuSLJ6OlZBKgVAbEmrL0zcCIfmfXXuAziJCpO
y9RhjKTbNL1LhX+AL/STGv5QLOwsso8yFFyjH4kVZNnD/9mipz7thVtRDcnBa8Je
GXgHFRYY94KqEs3Io7tCPwDu36bSsu0gTX1CzmZRv1n+4xuUEogK3/NWABNf9X+8
9jMfv9g7aD11B9VoRBZakmyG2tW1p1MnUvqNl1IGG2/c/x2g2EBgj7eQi9LD16Fd
4svCsf4EK4w/sJKXUnfzzg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
l5gMHgQ3AZJ4TzNQOcw3b9jawMQBMeeakJCI91mD0zDs60FCQ4rMjg0G/g830oVY
Sz13v07536QAi3s3HtJK2ub2C2B3MEkbsDt+c6Yg64x9X+VZhwvfW4Q6SH+gzF/8
jQRf2ff1KYlCBdwovc/C2hFve7D2DjQB1Hs3AndfO9k=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2592 )
`protect data_block
hSnY2ee2f6ZiB8UKVsNkMRDAw7uEDV274iNK7FoIti6jkfZ5zdHyUWPGxIvkutxz
VJwRLoMjP8VVuhbDXFJl3DUO0C0QifCJHxWL0FR2nxNwSiNKayrNuSPg5KdCr3S1
yosJMBMcpwFqUpq31e6oin3I+dEKLCCTc0xTseAEPARNejtxfw6F7/IBbB2FWBzl
574IGnxGgiSE92oRkoc8Cgda7UZMS4cpoaKHYACF82QclSX6G7BaGhJuo6tJdVvB
lFCoMbozf9BdqN/Omo9vt6vKvK772dQLXAFthcPBkbNr3SpscQpxJEXwXNWTsLa+
s1iJT3tcF3OrxTCzz1lt5WRjWWRMFLn8wdJzPIxpQ8MEB1RbuLL+R22dZpkHgx+z
rDLMONI1DlzolrG6B7Lpr6ObD9iC9FE3pJxdsyCPCUTkYNfCBimUXeUeEMfOSldT
gqvmN/wHGl9KydbmM4VcoTCfR9a5Vk3hfcCFAhy5bxcb/7tPjbZF+FoU87DCW5br
Gv00A1nt69PSJJKIehx1OGhJW+u4zTXqtQ3lIoBK4W+a8BkLyob82FrBqtiq0sxQ
wqOwsorZSVfTirRunm/VGNKwb29r47/uZ5h7n9bImXTn18chU/fINRRFvl6eLpw4
/8uqVZqpQzzw7vpVadp3bQDMt00X7Do4Qo8cAJ3dVvjmJrWIQo+aZxz5RpdPy8c5
J/+LB7m/5Nt83MSE2LqxO0Kyjwna/v9u0F2lqPYc8iccJVW+4tquHYnJwLZMSBg7
f6+x0FA9SnBU9IcuTKuYn/VOqRQYKYEq7Dusa/2htOaLSP/tXXFYSyfUOV8VlGpO
GGumeF0ExsGUN2XzuAD/na1wKAo6JrVLg5Wd2ferLGfboPvqCzk/3UBtAIDVCVWj
ffoVY63L58o4FW1qIrKQTxykTylx16aIOSM+Q638LW8y5BI2+yb3USTX9mvlD9Nq
llRl//OE+k7kSKAbrbOo2UxMIipN+wR+eHkz3KammQd3LbNDwxS0uf11XaegUsVb
LNoPLCq0EykuT4Ur3CdaJjUjqOuFo5JaCbpg1sWa71LAqUqAdW7sG6oIKPm8Fv4v
lhM9M/M1tXCPz6XAgu8xwX7O3tJvNVRnZudVqgLo9Z7nhaPELAZ0UrsaQwGzHkJa
cMAHkzyXljy5+mt8zuIalN5rUhZ7IpuVlD/Irek/DzLtf8bBPx0nK+te8a0YJVM/
3rYUfYyUdbK/PNZb6QViB+HorSGGUIWDewLhb5DxRdvTD2ZCq4Wdlz70Y6btTSp6
wQw0OhB0g4bpqQIzkMBxW6GXrab0XWioUxL4CkaJ6piyvh6Yzcu5GsYY77j4v4AY
23SQXWi86PRESqrLVv2ewAx1SxoA5kkSMDaK9/XaTCL4XCElq+PaiWtz+2BwbahQ
/BrMAwzRvyrSDG2nnlGg3bDEP8pQh1lcWr2H14cL7VgjPN0PrtTzch5f6KMsvxjU
zIGJUUGC/MvIjA1mtCZbQUAiXEWU+nFEhz2lrHDo8jkBtP/Aat9/QWSPUiSlTJ52
UhH6zKsIcaTAKUsrakuIZJiw4/c+hCm+EfEcULmn901GMf1JJXiqSLFAyI5bEnQW
E0a90Xmhop54a5lqP99CfVujyZvfB/OJexHfoWaUh0oHHAwrcPDZ+pLXfYlZQPVN
U8n1SFbO8/VBmunWetBqOKCSXAW6NE7KO34irYCRi15EIFoi1MB5TjFJ8HvBHjBg
0uWgw7FI+98XcjZoW+CmbO+dac3glLOMGHsH6Qc+2ry+fIT2QPQKlCQ0mH/IZ5Kh
OH4Jb26JYii9LIdPVUas6z2EpQCs2UaqhdO7YjRRUtxnmyFsPK0MrAz1ipaa2KQm
6VJzmzDOPdncVvWz4xib7YO0V7y5hINy1ZSUroge6rV2Kg3+dOWeqeufpQoWgR3e
5yy1gsVN9AUzwU5FNZ6QxehJDMMlzqsQB5jkuAaOM/G86YJypYm7zYBoLOTLnL0g
UBqD4mS8oaB7Q9SS8Kqj4MocaLrwva3GI3Dwgn39+e7/XA7DvCNbrdhepkZ0roAq
buE1R6HVLNUA0oxIpTHzf+sCS8gOncBFPBy2XxBo2P/JoFXhZqKL3vMOqRhgRjg9
dHnnpQr9Da3VoAxd4rh3FGX1UrEQNC+6/HP+E/ZMRaHHBI9Pk7iLzQPoLJSC42mX
qM0krvRLRU3ydKM2k4gYmOXCa2imIaRJntFVy853qvXSn4dgxrUEVs8oaIzfneAj
yyzRPKgMnIsmFwZYv+zrJ6nStkuVRioBZz8q/tUkYvo+yx00MnXlebl3x/F2FJB7
LDyVJILwLGnn1NfJX0QZe6mgxOyBObq4GXOV8YfN8Gbhxm0DESU51bX92wZF/S+M
Tj9HF4jpbRbdtXdmHsXjP5SqtrHJb2AtvXJX5eBUCsDjAk0guEjyXZ1Mc13OilRq
QVUzk8xD2uC//IMk+5K6W4NGWsGm/b5vaESIB7mGHvTPykanZsFYvN8WsQemYeQj
FYmVBBbqOrAZjNjVxWpEkH7X5h1i+Q/gtmiNc2LptX9s/c6RVqZx8EBGMck0svTA
GyIZqRkRkyoljCl4Gre4/VG1V72enV2Whlm+2anptHHDyJn6hqchasBfosY/6aPA
dCryh5RgHohyoPoCpVkQdiUHlFgH3lBG2/zoaBJ101nOhkkxjUUDy3wEbI72upkd
/EVkcB9bfaXxntQuw3ppa/t6ycW/zJhKcEIPcasH72Eq/d6dNHqlf09+UklbKucm
QF9qtWKX/Ee4tZDyfTVhk6T0YWKR31NMhyfsgeXcC7IFUpQUDKGMJVCIeisEbIst
pB5fskmMIewy/ihAG9kq0XA5Gx18Fwak03tW1bp87CrQZWDqAjHgN5O7aOLx+sGd
j2atAUdZ1d5e/hzRi1rZqzlWe0Ce1AXzoi6WF3Qktvv9COwKnSuSmt+/6h95WX8Z
Wd1lS4pHfa3bcscMMqCcTV2Tf6krP50R5rP/jlxEquhdI3bPjyTuz8nqSxpBma95
sW7626BfQaB/r8IMkf9kNWYpi1lgt4oSRXeyQ8sMm6D6vo/zLbQ9CmMZJaD4btKl
IM/Lamz49uBNJFXCaD1HspFQVt3xG1cy6pL5L/adt4p6UJLHlsYXYN5bT5RJLxcd
OrOkXDhAG1fONev7bR9RvwFElWMMphOomlHOPytnhHqvYSzTygBK7f55w+G4Rb1Z
BlbA3YTIemnndLse1IJjdpJeu5xgdN38ca2vueAPCkKoNk8/vw/kSWDQsWgbQt1U
O6pj9oUgLiuMtmmgu3m0NV1mkPXD2RlLtd9T4WqVSYRos2IMiLyaiQ1I3k/TjOEv
RqTFaE3HYG8zutWKuE8W8OgMPIte0J5bMQEjzMbLIQqOv3aVpp1pya4p1ljY+HAM
sjZXD3hhgIqfNirrNjwXwdxCi1LsEXx1LCMPIkpDfem4ysKQZPvbuEvBsWZOtk8Z
`protect end_protected
