`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bj5J/R0WJErJLOotP2NdeSEz7Q+r6+hVR5MD9oytnEtynLIFWLMDDOfSOyQiLCGf
DGNk10vYmKzHmUpFNf4LvjE2T4BIwlKv8q26KomC2d3xzJpzlYjb0ARvofZZQphm
2gPpmS3Pn4rEKERciVh9EH4uzMdvUnhxAvRqyXFb2zU0m47WiJadmrWCaef/YR09
P+iekgxdL+6Y7QaKm/DM1mDOu7oB7AzEbHEyvxuge3Ii0sANHdYjX832qjDli//C
pXsc2pnWV1FU0vC2uP3spWZL7VTe1XFLZ+QXv0sfwnFCYt2YaCUE9QdJPguVX5nQ
7gfnLunJw9jG39dWumOjJw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
tN6VqSpDJyIEopj44b9A9YSYtfCq2PXaBEAQ1ojF5MICbCi6UcddUib8Eahhb6HA
x4BjAhwUi+NKitYrruSD++qYHzn1K9jn15JX4zh2YaPnyYknd9LwnVVaY/RP2d7C
EMhqUjVpO9kyUeSoHjyq/UtPA//WxbIyB41lPDV8UjI=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4016 )
`protect data_block
hads240n9zJ9uldQss85S2T8I4r1Fft6A+Q5GCjldURAtFCBh1g9KbNljPlu0fxV
w3U1woNqve8o4+wVdDJSCjGtwBypqerVIhoEue9m5hSzK/o6ih2aJRhJHTmcsR9+
3rRX89Iy3vtG0F1LjgPsSpYCqhJbPp7bQxUimqSRVOgaUBE82hDQTWr/tiZNC8zn
ivdsoyrpav/86U2bPN6amiNi1rCunruI5WVNnIW+hJHYYVHKsXxLMFhKWVr7X44K
sw2WlWWFo5dIthZJj/quVoVouy0mRIrNl7C7qt8slRCF8t6VVKs7tAC3bSjqwrvF
l7Ljiyp0/nveQfEkhAsAhcYHT7Y1filR2iGqZY6NJfX+wpbkPl+d9ixyEjtKf4+c
WbL9LjPLq5iltDX9IS/5YQT751wVOh3Yobhi1hUji76Anw82cJOF9Q61LUyWJSVv
w6rK1miomehuO36DRsGx5MYzcMitPEONUuQwLDEgvCzCTJrqBfkhQ1qZ3/xPOCgD
+iJfa+P3PYYtH6Z32W7foKR4Rrcza8dI6VroVXDa/n+sxLPiuvq7NLGNArLBKt6b
zS6umXCR+6XP0yoTPHVWDOQc9olJ3VjejGD2vOKpRfC3S3izdRjkJfRazGlb1CCr
yxgC4Jwq+Qmoh/mdek+liRxw6qLIqcCVlz2ZZtIyLdwINfKefr6gaG0Q5RLBGrNi
Dbc4AliJBzdAPu0Fa59V0AxjYC1BSR+K4+DDi5IwSbKC1u64s/J4HnBvLK6Ndgez
KI6WJzycUXAH+w9hw3HMhpkL/ZKGHYHYcBoGcXBBCRUtPtJZmpSo0YFCvEXTWMjj
BGT4vZfyxSUhdxoUoO7y9Rs+Wkxuu0amTHaHIndPB0cDBzrQYqU6DLOPxAqGxcgG
ZeWqsTvucNYUT41naHHuz9+1vND3DrRyQMEskgdFDeQ9rTxQZpBaTMCfMiFlCHcz
o8iAHoP7mzev3WylwS18/9o92Qdfc1KAo5vbk6PdmirDHQGUAb7SYGL05mDN0Oz4
rcYd6VbqGWiPNRHAISVIUjpJBvDGuEbwC54aCwTi0zN+YOc1c5Efk43gLCrYkGrJ
y0LJZ1uxqnRl7GbvVzUdyMeajcPQyXX3DNFap8FVsyTBbsllgeBa6/5dtW3bP7Zu
kN7al/3f05gfgv567ij//vVvFN/tAXxNYYfEqV+8ZxdfTlTNqMeu8nl5Zzr5sHLa
eQ25f8hjZdk1tcZ5TUAuH7wOAidtcpP6k0RjWvV/k7eH5O+k2xcnmuoiRsnB1OFR
5bRADCvLTxdLr6pPJ2Ba1wpHi1hF9JxgZDKP481n5+SpTWgm63DB0SQrj/V3VB8u
MsdeXEElD3hTbrVz+K3uNm8W/y4s+HxP6Q21TjBj0bjaVHumjRVV3iMkrSVmMeN7
7BPahqOrUEziLmgyxrWNabsblO/fu8uzqbObEr01gMXSVtP3rqMSbKgK4y0vcw7S
67DC22jj5txyvlLehK51YNi2lEz0yGzG4oPZ19NpnZrrM4u/4DWmzgoelajdO53w
PKxfjgn+DDKO048rMcHO41/NRh9gEpy624RJliskHun/sFw0v+TuXvBRy8yjNpFo
V7KZaafKHUWCZ8+jblle+aECFsAyW56FImSXNDzHE6NPQdK3YlpQRUgwA6E5jQXS
G7hc0KpirJysLjRq9MZZOf2QEGJ70B169o+0L+JxTEZ2H3BCWOemdKFoy1oAXDRZ
A1jGFjnoQ0MaVN0TZVOf/ail013dbVmg0enePWO1vpvFJdzxW7Z/3fvsRHh4Ic9b
xtkJrLOMMszZVFa0N4KQpvNhEiwXh1ZD51i97642imaoQMpa08QDH8BiQSbJgu/O
navOwamq0n0fslmLZi4CdLP7LEtPuhpBDv7Qcc/OE9fuoo3Ljc+Knqma3wlhNLiu
SBnDZhkeyWNr4AX6L7UW73Ah+4g0l2sIpVrO3O5oXfAGegF0xx1qYi8Nb2bDCfpi
T2tm7ow8Al35yjPwWoCK0qub8Eb0Dutfa4AwDQL/TO+uELYXt94p5GIJwICELHmG
aBb+I3gcufnQyvxDVT50xpXZVrjOal1auwsR6Pvs6rE4yy7lMQO70xcjyW/sDgfG
JspXyTMQDyIrfoy7lqwvyA1LdRpG1IGwHZ8msn2QScsISmhwwEkU6Il7WjsmQptD
P6Mkpphl+xHpEUDdI5fcNQWnbHKoCvpjmKvQXRAmVkz8msHCsJ3uPe7ajS/ktFZb
OH8i4lNbIBaBChxJgV7r0+rqtS9GyAnh+X4G4V8N8C+sDrwdMkbVAHu5diCYVfYK
2iTD1OieX9NKKc7EPVj0DpfilfSZonXROksE7ijWQkbUv/N9UxQfJ+wcQTYXDDPi
Ue9ks4qhfcWyCITb8wUoIzuKETmMCtx4uLwgGGT+34c5TNWgSRxwPd4l5CYvHEqC
ZGDo3/q0cKDkKIZ7PGD6oLmMQKsuFscHWBonUfk0nVR2KixMY7yX77YL+Jd4dyg+
MvZqEpSkc/3rzxSf6U7pN5lL7+oK0rp9DZFOq5rACvITtQxgIU1kZM6IjHUL0paE
bf5m3niOt4s+b/CSMqj/qCs9E0ODMgDNTOGMFfvAiSSKKMNcP3oNLJpBb4FQRArA
l8y1pk+X5IT2I+/FGIfuabir327lbIKLyuP4BhxCFRjkrdt+MpSGORsqaNPlXFuv
6Za5Jucp4Xb298CaM9u+1JTP2QE1PWz86V2HQADoOwwgX6ICFnyjura47UQfAs6h
ulFDBkfI04KdK0YDZth93Jdb4PRaoCEcSZ0BdmceRd/HiL5B7zW6BOeqtd/QdZ3H
x+5E8w4lxpPJKND3+NDnaF1i3PIq9PQZxpPR5utEbVfmrr+bRB5O81LdGtWPXlg5
nmy0IIOTcvPmMzz2ZS1FZYLnva2Gh78PdZUhyVV09aBu6Ul5S7kWjTAIjrM753ZW
TXEYuPDED9A9g55y9QD+Mwl5GcY+Gvg3bc2w6rx6LNuCdql1k+vtS+Zf7XlY8vU1
GLiywDBAJiPbO1LOzs3a9s7LfhgH/+OFzz+lTz6zqz8Y5hH5x4SBvneKm+5KiKwd
yPV5enxYdFORpv6wdU0lvlCGd9hGVnbn5AaoHIdu0gqy8ex0mmpWLNH/ZeeL9Dt2
PdBSyDkNWnGlOOhYIepNYJOJAwf4eoPFY49oe4PGqOBi3LmY1CF2yOQNVy72CwJX
EryZvyACMOjexlcviF60dOzqUZb6+wypnS7BOW67scesZu+aCwH7m8El87qreD70
qEyZJW5T+VfOllE8wjHk5AVLzvyrrzcZhNBjuR/5IlkqP7OTTCwYD0ywfc1tFCjf
mU9iU+qp1rUGr1uIot/ynTDV9vqLaOd+bJIh6d2SPnjbq2IhgEQpgrCnxCB986op
b79VvJnrrCp4eNGXM5R0J2w1n120ig/Y8ecXy3PX01ye2/ra9gfbpEK97J5OEO5t
nBh9bqgOioBK3u+gpaX7euwHlguUFKSqUkhcj3j+dwk4qG37YrOO5t/xwWsN3UtJ
GvsCQQx+FNVA40JLN3T2mbbVttg0AIPVomP1DPGkcgNXCAfjcooSCeJOWiaCy8Dw
dVxz4ZVdmWLYa/fCKpQXcKvpAbib32FOI4Mf0z/jOjCRTNdPFNwUIqGBbthcWWKZ
B0Qi2FpzeB6nZnTn0NfUwitLckU92wOC0VXHkl6ZQDl1zmcR7Fwqh8huPktAk8mB
YrSppeehkotj3xC2vrDYopYt+YL90TCMeVyxS0Gy/6d1CUTM/AmQziW9OeQ6ralE
igIrZEyHHcH9Se0HUvgabjTUQlauSj7Zbf5kRvJS4p4AtTGMGmO0z51baPKwjaJg
Yf93UF4qCb0f1qCFgbBWC3sCwYc5Tp9MzIa8nhSvPST34fLPEjO7ZqTRaaWdOsFp
oqrdXfPmT21eA0lWQBgwkliMAzo0bjHv20osHnZRTk8KBISb7hrEC5OqWApwFJDf
BoIWZzSNtd66s7vVHsZHFQnu+9WAzHMJ8a2gy1KrCt0ScnsmUnkb2QDQKcuvLRFF
wiqg3mP9Lfm58K+LQY9YIRVc0m6TkqVd8IhY4GHZP38Gzs56yEl5UMoPGaO/U5BI
Ao9o6bogUO/MziX+WE0YPlkWX9idu28tixfG8VEOud6TPrGh7KkIIol24XGk0bBQ
53Xe6HIFdfZXKcJiMMP3VqJ2GithKLOREsg61Uj5tJHKlU4TyixVs1tezK+Svmv6
KWGs5bF1dV5kkHPtKZrbanCwhIb++L9OHKRNRKJyOMsh3B9L9B+c3di66b+FKZBb
XQPMoUF6YjE6L/hoF8sVYe1DWJ/ocBhQyCCRjl9JzpOfw3oebI28dIdj0MI9bSi2
gbAx8wY/O69mam7Yl7knY3m2qicZk4t9xBBqAvP2BPMSYFquh7n3dU+tJR7Xfv53
5iR3LmHfhGM0lBA1YToj9hkGB0/mqkVKC9HSBTBR6DWHWyTIWVYWAagpXZMcCDf7
4eAFE7fyIejSQYp156kIg3pZZEHZe2HSGGMxBdylvJGU++IdEpc9aFl6TRn97hA4
r5mvzUaf3/7kPbBnNDrZWXvA94APaJDQGejL83aFOTt/LGVRgBIG9vp6bLT4cFYB
+ch7pYLB9HTenYW6245+aZNRl3kEEj+wPfZCux7UCDKnY45lXwwB6meGWjXjfZvw
NZPKgUbjgcch8L2QolE0D0QAHdnDf0jOUiOB73S033DvrSsyU/H88voQxxHHwSfe
w+CfpxpnJGUiuKDyyOm98gvEZJk6AIXKdbCYCCrFkF/d0v6if5ArJyNUvxNj+tln
IZ3VjKnZAReTVvB6hiwmybiDa/K2ar5Oz91DKumOe/C78hFgffcBNeEs/xv9ZASH
5tzmJ6cT951hIta92+yb1t+TA+63Xc/RGu/rsEz2CgHha7va56ADoctkH+MtiYS9
s1a9Og4yuHCcp4SvJDyimc14N5Bila8ox0GdX5agskoBjkFemorf/Jeng2HQMT3r
xk/sv2UmKmlhXbGfx9DorX77kPH7IvzphTozqjYunb99yGWiV6yJ0rlvIOSAuzfd
z29V38r1S6R9P20Gz9MlSD3OvaLdn+Utahd0af8exJOtKiW7AbdWfriRuuQH94eH
AnfSmpJw14E87rjdepMye1C1SiEvoBblTRXVRUGuoBrnTbUXj2La5fWcuql1F+Um
JYODJ9rVSF1NkvcrcnS0BAtznauE9w8uhC+p4ZFZgS+gJkeGcmBiL35IyRELLApj
Rf6tGjBNaUccmEXllo56HfEVZrzMZzqow7YzhUetuyoAmKe5ynVSFQKzjK42QyWR
Ytd7InWbBsrSxb5Bl7JrdG5Sd3TH6iS2NoyzkdkNSng=
`protect end_protected
