`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Ag5y7ryKz2TUC/JChUuk8PJa6x7xT6v2q/GaMM6dot/FO+ChemZxR+GGbRT8u/GF
kP2k76fNM+hxydCPZjt7LA/bh1iPjAAAWJhV9eh9wDXEhEc5wT1lzepdBonWH/B2
xBPwBW73PKnq3D24Oen7VoJgFHZzvxbu06DnUXfHMAVNnFLhxrcDZE1IMN580c4N
/kfoPABQtphElVyCuVm6cVqkRt0dmPP+QoFqqLryzJnqrlycFWaZs4KZIM+QAWwE
sJxxpdKkIaB/Jt9rvN0W1twBMw1QKxcEeRNkpc7GHz/nKJr5ofo6enrcahZZhcN8
LLP9QuW/ZULMQWt13xYJ1Q==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
VmVWkOkxVOrpxi6kN0xlNOngnwMqr+er9A0T1VZKsMQR1iTmqKn+CxNWYlK3panT
4VsKKpCfdoHqGkChIn1lQ5GDMIGmUsKLk4XuSuajx9P5/sgbwSJTkgwa29JM1Wvz
kl8e8TX2+SB/2tFNCoggGDVoBGAo2KVW2OPOgEQbzlc=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6912 )
`protect data_block
EfDPrktZYx3y6oa6+WVWI0twHmFpcRq+fbB1IYCRppLuwN0smYdm9O9B10QMtC9f
UJ1+jwE5EiBYFbLaWPhh7xIzCf4tgARSZtkdU98NmIohvi+RATfpj8zGFHOh3WQA
DjwOewAPUBX7zzxtkXfCAFmxAaoeybT3YVl3f7807SgjugOM3YVG86eGRW1R+ZIO
sN6QLOtDurVNNWvQrUL+jTSuSkIxZbdXd+kN86SvmRRCUuZwwb6TNlgb9LeDIu5f
6vYrTtaXtO4GgYsmoRJ4ejgrqb0mZ8tDebVAR2AdojUotR6l2I2yt2GEAGhK02Ra
rraaJHBZoQ3VouX2GB9ZN6Wq/dRuMvFVhUagzh4q7ED6H5oKYvIN1ASqsXcXkwGn
Uxvj3Ysxj5CG8qbl5xgj0IyxA9xnb0p4aUlHtme3LuET4jwTmm2z4ZAZaPyqILRo
fEUFjn9lkX0rEoYQipK/dc96gZQxROS1LfN/fcKJ9fPJG282RRKiN6YSVeNdHgxD
XybnZjZ2yLHMyPsfSb7rLpyKlmS4rX3fUjzXpmDVpwLaSu+fRIvfT0Db6yIhk/mA
JRG/gQMEM6YlRmpu4R80t4k87FcbDWJoDtTbis7TgLz3doT/DGSEoghgIlo+Aawg
v8sKdcA7Ki262sSFsXmzCRHQ1wqTBQzYb/DgOfoujxPmkJ5dSSpz3Umf8ZeEy/yH
IsTjGYdhBe90VkpmylLFvhlz2EXd5kgPe23KR3n2VqME1adzBFZwZPdiXscpvBvm
JbbzRfAuYuNt3P7lgM46RCur7gQqItmbNugmR46mICKPq0w4J5+ygbWWeMMhnf01
7NK59d85Axaogam8XFdBc9cveDdkkHmoRPiFZz3pVumhm1JP/j0Hr3jppje4PgX4
JAz3DrkQ6Oz4cMXo8ZiHr2mrHOoWMaYJYhXtqPYd5Q/eeeS0REeV0biqn7KSPhtL
u3LCD2PMgdVW4D1XnoU5X9DK386on2oZRzYnhx4soKCFf0/Mit5XCpEiH15TGl1J
BFoQFdgpgY3OL7SJu66MvFAgQnKYpiA1b3D/kUZ9gtoIbYtzcvp30MOmhszku7pr
ndzQnjbfKTk8eD7W/F/DDzM1p9zTQQWUIfEj1kBgdQm5gS5ER/4fBjdsoCF00sSC
CzY+EwZn5Y1ezM1v+Xmfookt2glgHa3QwoY15C+Usk89gJTxAWJQR+7GRGGC4bCN
kOAxJ6oyPvux+TjCZecTuwRLLZG5NKeGCb7pgi+YAoj8UnQeLcQu9Ys9Qb9WH0Je
gsmspbjuvT9WmKVmxkmfSuX7fLiiAJJ1j1YE4vEa5QU1En+tv0XgdRwF1NHlV6Kj
iw3yvhkSlc6D9NITZ9OA+tGZw04HfRzXUR+Jtg47/usc2j8IRE1TpsBkFdxh6Txc
gLONUUAVr00JxrcNMMNfnzDSHvaL9A65X0LZBGS1GMG4r739ZyWCf3h9hghMIJsJ
XPEkroJ2Hyj4UX9pxTGTObWBu+nQTb1Mq0ZgcQlZCpV8qsioVgD8A2Ny2Koovkt8
y7VYz8joY8MxSDrlSzxEaa2hgsnwWYxHJ1t4ypMO4YXO6CRD8+dSl3l1HCAnnRoR
SgbvIC02xueGiALlNjiepuGBFnv6PNKXep4R8kwxq/0rEIBJnJ5bQWEc7JLVVh52
9Vo5N4gf7by89KuHfh4UTL+9xLZAhHvntSUNsvsbUac5ID0RFuoejBq2WZWclYX0
Y1TFplusOoQ70Z8YhPcC+Qov6oOA69bumbL7u/2NbNK8B+i9JqLhaUlMGKkGkbdb
FwqBF8I907sBxf6hUCGQxfx4CY+OgVNFaORTy7RnDOo9LvphoFq+7YVQ46aZG588
NuZzbPDVWEX8M97cww/I+AWA/9LDnFJFrHxuWkMRLONZk7KJ5lxVVg8ML8NpX9hn
h+XEbr8v3oZxJSjBzE7jKjRhpgKf3rOsmVhZyollAtD/k+CIy+cgO6xsAp+qT5ka
028h2ft90O57/josvetATcuaKIL0s56600unrSNfSRfEvFGxQzVO9MKrbX85vFZy
VUN0J0BHsu+Qg05kMYyBwvGzIaVKOZeqTYDxJkXArxJfAC1dGihxVWnUftQzMsrf
j20gpr8iDXfw8d9jNfOdC7oUpqtSeKyhXbuwVqzdESvtCMW2ofnV6n8cvbdkx3Cc
avH7V7o5efjmhImHx4yTAgpGWEoC2Re9VNvj7c7ML0m2PdJZslHO97RENdyeXpeZ
Ejp16fRa8Ol9HeSMP7SbZU0t1GCGUvkIv5xdSi5OgWsm4Xv9jkt9cGhstG62SplX
ZxHtdXbgNFDGyjRjF8K579I3D9lGXr6yGkmLfG2kH98iKDVHOzC+whePfpNTkIYc
QSLBjzgoAFviDrZeiTClOwkfSKN21oAjF9Pl11pa3+ec9MOIBbiXup7cKc1fB0MK
a1AsRHrPJQNFSQ1aK7qr3kOiU/NeTnieWPoqGhZAydtNjm9eUd705tdWvZeL4Bgu
8yzXzFyEh1fpzIQUs0c3i7GerX5Xck4NP2/s3NdoDwcDm/I09Fz/CKz6MJc2oCfC
JKGZQm6jp/RGhZu9pBzv9Es8oqNGDroaMVVR5c+d/aY7Mh7rz5ELn/gUhYAHV/YP
WR0lR7gsfTKCHTLMUaiKiJAi5TOkOhdtdpzggWXwFW+bUTfNUli6bl6dM5H8f2nx
BMA4rGQydmzmMQ8iS9y2OHZl1esHH2bEec10ymmdgXh8yhMOlK/7XeA38DEAVKXV
WyXljBG0jwF0q2hY9cPBa0biJpkMk89qCbXV6pHmH1I5KP4AxldkGd7MeYEByU6Y
6ivBR1wGpsFX2SAbavH+HYqRJh40afCq5GoIhhp23UgxRXEEtr5dEqz5P1DZQNLk
w6mppOwsygurKEWF+SJrTfAsEFwdkMGJe01t5BdrTVdLo9rvFR3ObAlr2rka1/yL
4bB1aH1e2nwEazW6DxaeaoGE4+nASLICXs1D56Wc256Sdz/Kads1MJfEvWHlWHTg
a6pXKnL0q0M3to5FtIrelvIqHCTC3fBg7G5O4hG1EOq2ripf6aY6EgBIUJ7wPFjz
d08YuosZCiMTLrZ+f97deGK8h3tl4luwsRmKwKYNJ7i3UXwg2tWuh59zeBoidX4g
zDREZTEl3u6adBID26Oz9nw9vedhQx+XmJrNKjxa+A/hSnXEaKkMHSrE51EwSNL4
VEXQ7iMnhhHFu68OtNbJiomYAVLUXjm3XvvplEglRDAzFrcnNHhH0ZzR/5qdNHun
EDlza3JVM5FpVP/Jw/bnNeRfgPvWrYx5bkf457OekdLQ6UUc0meOZX2GzDt7/HbP
UbkZHUfD5fBd+pFoANan/AML6oN9NSwVrZ862eP1qdwdWeQODfZIaxVTift3rHle
kgYLI6nU5KCqrgGqSHA0Q0t7OSgsd4XH2x99RL2LetcASA9lUDBT0UkkIrOk9Rxs
y5xtA6FTmn7ieAxmD/QXZD0Ba6nJym69cyGkx4eTER0Dbctk8A68VjLw2Zy+CLWY
2Oy0ahs0GajB+Wz4v1EcsQed/QDQZfRLNXKnpjGtiztnWE0EqwunR1ty4lCuTEFG
9jA4/x3eZ2r2J0MzY8Fa1fgpKe+NjQ0mE2U/o79P2zOmI4ObM71xQbaOM05Upr/4
Cgyvlz+53Zv22l5WwuGISy8wudFNJve35RP74EjnR63DpIZt3G/6GWsyfJMp/F3E
vu3Yml6gko4y1Yu1rUya24yf4UVN0tURokSpzhPkJfAXr36FwvGgfO6prjT/Y6DI
FblXqlsPbSFwC8vfoq/Xd2k+AiK8Pk04vfiQo6Zp5+hR27DkhYeMSxrS9Ym3YuYg
z+sOlv1jy9Ps8nrnQwCfh1Z6lCI/x+wXoj76tz5iLYtTQywYFXDSYaI4sVQqk/kS
1Cxeib7c8sGq5CyMTTzJoQx4Uw4GxxYwvkVrPPNWFZE3AzKSznYyxTHTaQqh3/eM
qmmMyEGuOh2kEOPe1WQKvqKN8xM5/1LFeLDwzl3e8PBtiWfuVRkzfCHJrgOOf6Yy
yLYqzyZ6kj+Mo7Pm0P9CoITJbs6+E/FIdUa+x9gx+OyPC376BUs1Yi8pKmCsrErn
OYYsMP5imfK7wHc3K+1YZXKgDLI6DjzOB+3ul2Lr2TXgh+N+bzt+nxtNXUF7n2qG
Dz/2kjuD/dn+n+H1hbXs+Aw8fGyMBRJls8artr2dyjfIqHAKKlzvOGeDZzqTSYaj
L7QfjDHyzOdprWAR2+oKTO1JqBHvSgFWgrOR9u6QSskAP00H2mQYuUL6Ix1nL5Wt
ZBdl7GrkwlHdryAUW9xFdC3uSqct4sNCWZM0dElaA84W3ntGTIxWs8HXluBUXM2Y
8vELtCx52t2XdG1zlZ4o1K/q6ThvJdlhilb2ZAUwgAVF29yHbjOZwmhSammUBPa9
ZwbXhagQrFX1TojNiz7iLLFqBKvroyz3O4GlT4HyUzNOvC7Cbqr3PBI9eNy+Et4f
m8yMc47OUoAfzGFgtbMIDZfV5vAQua9bD2s7TdAkp4jpy9QQN5a+YiLzx5drsALc
COLrqCaqOxPT095sqJq+JrhONqsqjct9Ie/cQ748wHm6jCS9deDMR6WxIZP19DRI
7PXmIVs7H3DsLPW/O9HslE2UNbS/pQFFsKWxHGKEDmuRc8dbdyy3QTJE7Z4MNBro
DoTSuxkp7V36YWqv7ZO7QE07oFysvDFVnlOFF8hAScs8t1kTa2gV7LG5GVFfKPVw
ywEa4pkX6n88eXRDeSmkJxYDm0COgG3zOVRckImlLXXcV7arN9a3yTY3Ty0Rcwp4
qz0uXNcDXty1liekpWkUYzN0C2phRJ8g94AQoY+tAJbPubDnYUZCq++r+yYJpAzS
SXvnkDWa1D3Dh1LmU9bwPoAhQGXog5VHp3sNUnLuG2OGGjUbLaQ4sb1Z+tnkVjhj
YM+axc+xd1lDOeGKKfuBHJ2EGUI8oJF+BZqg6ao9gz6Cg0K5SETAsD2fVWIUCT0J
OuabBwYt+jjazXGzSlNvbkOVHkZsxMlkcn1qOTv2Ng5neGhhrxpG5/bb9ykniL3n
sMA3B3PBsOZ5f0bek155Tvcx0YFEARrUg4m65RLkwcp8pGbkDZhO2YT4VHmZUPfp
/SmTCM4YmayTpNmzVtSEvncj3nfPuHCqF45SWHWP28nrafCYGq6q//b3orMp8RkQ
R2hPo7AHZEFE77fyr5H0x4vKjiCvM7Lpa7Y0vqMQn0RMSanSXj7huhEuOLyHfpTj
4C2tNJ47isaMqoBHY6APUfhg1MRo/Iv9/5WRDkxms26nbKPy2UABDseLJJmThJXn
rnSPMkUHtAdVSUwsh2nzct2d+bLM4RKTxeNfcgtd0pRXw20lnFneslBsFF1boWWe
Dy6qIm6T03Gye8ooLmwoNdhznCaGmoP90jzPQJ0emiYGDsCX9mL0OuHqEXFVLWTI
wZQG/q3La7KUWA8MIXZyqYaPWrc8e5zLbg1Xjn2ZoIielj0VfPmx5ABgYZB+GpsQ
FP5TlYpyRNxuS24/lubCtgs9LeupBMFDOEJNG9Y4FaootKBwxXLoRAVFh0bk6IbU
haMkn2UhKXJjQePw013UoRLOdUJekrkJS8n6NlpqUyUnxqXRk6SEGRzzlrQNoaMe
SyLL1Er3bzHY9Hfijd+0ad4c7YBRd3vNzDLDqTdojbD/OwkUrnro3ImnHTHUTcKc
S+0QpUNMwc8bw0EweB/0sWMNyGvElMj5KVbqTT/I9DNoDrNATGnc1LrBWnB2Gb+i
9sOvZd8zhkx1BxyzpALnfMlevPF1OdiSgULVntGDVZrVnQVZmABp32JwIBQS4lhO
ub2fNivZij9nDJzxb0qTTPQXWWiVLt9B4f2Py48DTAA/6dKOo6wWJVVeSSjJcwZm
+YfBbSRkNLkhLQGT+lxRdOk9A6yUDyAeoalg//6+TF7a+S7gT7nhNGeZEDpDuyxC
Xxg8sHlpDPPpeIoqBAJrOPp1kZ8Q6gr5/AX3XjFACT95hV5X0f3RAtkZRYRLIR7G
FuC+YEwyxtYoggjYCMP9mLuv5NkpQIfIOPoppgRq4pfgSFu7inSvrZJIUw5L8bSN
GoeXuL9uDiR+hLm5ldYQNxFhUE5ZbNuwPUtMAQnJbR1bugGIv5/OQCiiDAs8LCYk
Wtkdb3sujxHkwg6NXvKljD+NLKeYuAvulKx2ObOu5w1QFwSps/oXEwI2BQUHsod1
pONI5b8zwe7BsNEsl/cUorZVmtZljeAM2j3HB6VYfML1uiF99rS9DhWNesrsSchM
TG+MUrWyfR4BN7a3vk1DOTuSx49azAzSx/5Vq/e2ccWkwuPKYCo+aSAzaVagzP07
CfvP/VzpCPok2EobzCcJYMYpKwyodTOPv8IMqL7y+x1Z+SNZ5bAyBUdylRiZu4qT
aL4+5UClmn86la0zjpyAmFG5cL+b713UFmoijNm+sPkOfDgwH9Ii2heLlPX2mFAN
acm+uiqiA1jjwyKruk5ebm01U3ymHi5Yzvn/fadM5ZlsFTKauItT7TgRd6uwYic4
QsOuidadZN8K0Z8gRMCBI3EBYFIX95i9g4kEokER4dpGnT28PHAwMeB781D5f3db
yCtNjPUcpH1m+ebv3AhlA21smC44Pfy4Mpiw3D3S4U63InIzNjxDVFAfkzFwMG/5
w0koFIPuE464XvvJTEXqHJLFvFrSdnTaLsFzAnk+alF+qmCUMK3/nHiUkzimgPl8
LKlG99KFxn6jWBK58QHat7x1cEwY/R5zpTOcsNVA2GhgXCUgyIofPjN6ZvfC5r+d
dPg2F9xx6VLZcoJFmhrM2NR/jqHK/C0sAQox49pPmRzdavA1okX3RJv2guABO3nj
cio5UX3E5T0y7St1/z5B96SqCdfcOel1zg0z5qibXI8kYxHxHWsO9DjUKOghG6GO
gVpI7tI6rMEr3/Yz4GgLLtQfWCLl87Vdt/dMgrd0NsJEnOuypPGZzGcKCG0opUdy
LmYHAeL52CZFP5BeYym5vLg3rvQXcd6nuhS0nNTD69JbbqEIruO59gtkoSTu16vV
BjEzm0Ni4kbCKKbsHSEkejgRTjfv1F20okCQuJ0yujH6DWQEzcD1hcsCcfw+FuRU
ptV0+LS4JmCZLFbo6SSFIyQUzYvoY+R+sJMjs2tyyz0Y34IxVfZANvv43GGouCb1
Hz9FNDlJFtH4xF4xGVdyE2ibiLtKKf/JMzOJFz7e1JylO2DB8u6iAZ5tlb2rus9H
1qXH/IbezGIlonD8juTdwgJ1owl7pzr1FMQB0U0gqAYCL67sttyFlmpQ0JJedPhM
z1rI0XXXnPmUE4OSKDuTEmcS2wFvAy3AF++w3+g+EgtfGzDv0hvuawittV8M6xQP
26gs+lSlFol08HVXTD+xMEtUnbf+qiorWbD5icz43vr3+zyaU1T0Lsq7nsBokmmN
Vb4ZyC/kvLG/od8k5fr7U7KVLTPJas0HJIlcXgYcBdNLfECtEqNzaQQ1y8eZ9Oza
J3w3KQAij+/qwVNsoeS8RrfFQHrW2ZhUrgH0vu0vvWAywwc1ABl00BbLpUZrtW0n
ofK4A2fxJzavH80dnkLiA9Rs9UcymDtoaN2YB/i7xD2Dd/7Q7N30EC7yGxRHS9nw
KYkxP7Rbev/ZVsW4Qt3vVUU+7m+hRYV6s8rWjp3RTZM0Ch8uNQ+SaQOWInYEJ30U
bprXFAuR5BG1TDLWx2te+QHoMsVazDlFoupYcD8SqoaFtjCYWdI2n08rX0v0tNVV
6JVhSaCwZmpqRgM/ntLRqvRx1DA28Kk1EozvGB5EcpI/073d3MaNFuusgAJtcpgC
sQBx6fGM0/069gotAjLhJJdFHa94vo0DeUmpw0VOuAc85ehvimVa9a1iybARnYu9
3+7JKXt8Nxzn7PUkYHD86J6FSJQzPp0KvJnj0hMFbG0WJdougPKlL1pAKglyA5o1
ir9ME45erOmw0uKXlKIRFKLOcPlXxpp+/HifJYm0btM0bO9EHuBzsFzxv1z+MW65
XExOJvwQF1r357Gh8WYLsgMFmRh01e0W9qCaDAuJ0XztkOQAOFQ7YyNYeQOaSdZb
kAtyI1HNTHO+dxLX/fmMRNbuc7YeOjHKAajY5foITxC5g7bhETGyVsjiImNCdFPc
k5MKDvTdicOz87m9fB+HAd3tZ2UU4scu09pfgeZXY4jTXWy8P3CIh0nZRH422Rzo
BXgHpsbwK6RMoDgRIX0lwis1ROx/h3O7Rgy7ZDn6goqccb6sNisVk7RR2M7LSARh
hguGJ217h3hxv6jtr2LyhBIREG4AgbXb237H0ilkJh7UTP57wnvn7rmaFLjbvypD
4oq+DmKUV25qnaP2zgdBE2Nbw8goAKOSrPWRuFoqRsY3ULZ5b1tdDO9qwwEoEtgR
kMy/uMvQByydm20Tkejil8nbcGFF5ujuqPBh9TWT30hYx+diySSGz/XO5FezmB4G
pNlZd2SMzWyfdf0rmoWm2ji6MA3Ue1gRzuJUpoTxm6qph0jZadqeVHK1Upjf3xVD
5jyITYJ64qDpwZ0HkFftMcNd4w3CPdtw/boF3Wg2iYxB7nKYo1culiHk5lDQMyzi
iInPIONs+jvIDOzy9aFCYw3c35W+aIBsIiv7QN8lErppjG1TPFd76g5GJ9Rlxvzj
MviVqY6I7thgICNl9mAQXZcmBdNcXxiY58Ux0UkMMYTJy5jwFQr1YsUn9RlyXa+Y
SsmZwVmDhp6J8/p1+658IPETJxAXzB6o9jRsiVZ/osR86nx8o6Z8luFb2h1OMjBE
bx/qiCC1zZZpkAiEv0cAy2pw+cpDbWpxeXjGh11+BCem8kk1wsiikmrZ2Uw4K3as
Zw2jek9WeA227x2WioxTyIJmS7CWmAUn1u7T1Z6zo4oPxlbqF+HXBGUcydymzKKv
dp3ORymidrgIa5C9j0t4BDeI14d1nCY+9L0kddNJXqWYqETz8LEV6GkCAN5J/M61
Vh7D13qxI3Kpbloq+AX4XpUVfWW/NoFeEUKvmPD06/Kvds77l94Pc+ISWD6tdBQq
HCu9cQYz/YsyAaPQBzpYmwbSeRGy16eL6GtmmOQSYqkEv9z0HptfipqSLWcxVJcI
Q+ykaD7AASYT71imLztasULH0BbvNZKCe6x42Uj7zg4y8OahfnqNwykvhdEuLaQo
dsUXnQy7fW+gONcjCQ4COsDy0GsyWA6cMlaBxFSzet+tclLyL7g2azPwg+9B8cHf
`protect end_protected
