`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
A2lukishtW6qBROyTFcl/pg+Le3EhiTS1PE5gxcrGELE6LdDxyf1TuBEkj+0XzTN
T/AN3IfkJQLrx7gvb53FujcXTVIijxzJU0AlWaQyg1izox5JbPwRrfmcLuwPEhq3
jfNWdBUWtmSg5SxwlGeEMrhK5zxwaFjQqO9bTOUiNVywQa6F49K6I/UWiY1u/xcd
bAGZaXNIwvTLk/q3exGndUNcU8POdIgvkeg78oItsx+RKOijqZQOUtsXmCB6YoZ/
K/A7PCHEwPQrnXKhbgIgQJ7ztdvVMAWGxMBRnx+TmTLn9tJuCcxUAJV2RynBnODr
PR4qaBaN69Vj8t+ogy3wTA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
q+BlYbeu+vI5FPcYrOnvaygPGMtvqWEcHIpCjtF6UmIK4YFkvcLTJg63uNQ7a+HB
aVjpSlMlN4l+VWj8mU2NrRfhTSFdxV/u3eiO12WpX35KJSMCQlNirdVFo1u3/ziz
U27iv+aECCQP2/1gojnYEqWjsi91io2z5UQUxCYA8l8=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5872 )
`protect data_block
wtNL2tdM0QHhd59M2rJELIlhOCXjkelrdsvez8AylE6wq6voQG1531CjV2Kx52EP
R+B8HqeBsPPJoMdx6HfNuTnD97XL4XslBsAtxcoJk39dOCZXQgdz6+WqH3B2Zc8h
UDCWgdqZokj8asnV7btgKRGS5TVrNuiQKbWsu4HzNB5ZAU/14SH/GiOVh8apvveF
+plSomdBIGsGaL4Pb27br88Av/9YUba7sn/zieQcOa8gKbRUSrkcgWYR+Db0fEKP
6nUX11A6Zwk9ngqdy7wdyJ99jwT2ZmwITldJK3NSSZ+VJvrff24F1AzecfDLaUFw
XpcQsom485FGSY0oyFEQyt0mYao3IPdowRqlsSkfidMJRdey6K+z7xwwQ4R9lBsV
KiYhi8LOwF2SY059zuiIUu8GM39ou7oU1IyqMNVZccJS6iWogeNGlDA9pW9of9wP
EYas6UMeC4O4oTuGLWev8teGz1mEW+ONBrryAZOnDRy16uq2ZVv1Z5+5y2dl8R94
UuwAHaoJ0/AgZHLrIKOBJRc6FD+3v6zO0RTo6+LrgxX8HvK5BUYwx/UwP5DVTjkA
eHwJQZzKiq6uT2GiRkuaheTGtdjlPysMZDJf0hA0zsvcFnRVNVFuKqbq77IDtBnA
1uFYJGpvDoPyOvAeG9tyPy/t0nL4xi564UFUZ9FYO7tfmMHlVaQrG3sSkp32EyOz
2Urdxeh9WGGwisVQao4WGf8yEKBrAygqMYA/VAfZOxRxMwa4yq/lgt72mvCNn5Cl
uEw94jQN0JP1CEOvQHUy3NODg44buaE/DyWhIa8klzyynJzYJ1P/RG5axzyZuLqm
G5OlhWrkdiVrVRRJx3+qTw5JV4hJD0BIfhR7NzVJ/cF7fdUcKGZtYcHVZsF+WjxC
kDlzHT9xF2LAyEI2CXjlr+rDtE0yFknB7fucwOmOxr9B1zvmlnna1X/1mrdOM13O
lGinWhvnyqhLIDJFwl5pyXCN7+OM5Nvnn8dPWMI+XTP+GIXOjUz9J74xK8KUxzwF
OOa4ggUVwsDim8GqSeDHFSVW4GsmyHgGc0YFfmqxzx16zIMj0PMpijP/Hg6QVi86
J5Ghl2B3tb1F02VJCV1HDOnS/MKM3YMStVVpGzF8S7Xp8aH59C8CUVQiwaCykPLw
OBVfuvmc/DjdL6cnoH6fA628OK4AzfPQmgTFyLsl3p63UaCQhV6UMaiCaN4ywG7c
lr80BWttElMxr4puTocHhXEouiMWphp4igz+bzOWPZOB8yA9gBqi1EthBU/BPkUd
c6MRbAIprElECymPlc9h2eD3yzTrXUCQLuN989jGaqHtZ6pAFKCw9j6N3p0AIjgs
02TgwBAtOyA9WCRaWvR8tfEkDXi/Lt+++x7WHXpOimqCkecL1g03hah8G7UgQ52q
4HnSBtls8XB1XPEVrrwpqYNh92q2zdrHiSbPQqZ1FvlN2/pR5A6C+jFwUx7136wJ
X1fgrRW2Kf3iOipqMP6TuPrl+/l1KOzJzK59kXuLZbrhNejOTk7uSXDO74W3f96T
rA374VWtyDtuoDyncVwRBwWssqc2E/ngue1NDnPrwUYRBtciVLcN8sIQ/3yTJt7e
IvjSGQI0E+jH3aU35SBfOaVAmpeMOWwJ6zUYQmmKc5c76zKoy+cxhQK4qw5mdGUW
x9FDoy46dOdjO68dTj+XWDa2pAtPaMlOSiHlfeSedYV1pz8YFGO1SLPRw3zwVvZr
s+VECtT2esPDIXsQK6q3PDAcH+PL5zF1CuGvpPv6jpgX8ek12zl6IEod+bJEhYMN
fudvYKu4G2gaEnlkkPnPAyMNzKGzjK0aNnazZXu9q/FIKS0wjPVGdAq+XyKfTJjj
3UdnhykQiLb/pfVLYneryG9enYvdHTOwcsDXMlO0NUWib3pc96vSHm1yssbzaGK/
iAzfw8cIFTsDCHDbJlqXVgxgjnp3XOkVe+l3PzgAMUGaJf5TMhZKA/1X0o5OT9cL
ygK03MdGVttfC5FZMci4ry3bzlxx+twDy6DYbp1I8ZSeRkZABHmsDjSJAtYwOjqq
Kf1pdMpEYQtWbXyghCK1UxnN9u4o/XZVgeJ4wvOgAZOvsJYqy/Q6xGoeomsQVhaK
/lsOb7u2jexGQm4nGksgMUPok4OeoTU56jzXI/2fsVyVGIwfx/NM/O65n7zQDIqm
wJVKkHmHEqOA4t+sU8bjOQuWdDNm56Zy4eSyUTWcj318WQaMPYQIyBlHT4EmlKSZ
NWWX7hzC0rhaBuWq0oo5mb91jdH+ZSw6R/V0Amyud/lmXENOU+5ND8wj+kwySJc0
4Tf6Lu5J8pg/f+mhzfK8YG0dZMHOXIZEllaxnsh+JBKo7lrLOiYkuR8t9FDSwEOF
wWXPorvZIohw275DDOpgGOIaZONO/cxIxhqeK98xlEiHeiDS6Jx1Exu1r8p5q+eO
AohbZCORfSRmJ6snLuN+vPCQtT9Ft5SDqXH3D/ig8QUySUgaAQ+rRwGyROC01Rzl
jlKaRKQ/cwzxVGQMG7on8WmNf9qBI/Sh/7Cpz6SYm4cPicfGy8j/X2maPZpaJl4y
g15Ii4iKzlkSvusJMPofLipwr1B/X9xhnru4ZibgGL82KfgL9igV5h1b9DuRSsjE
DyfuMlS/OwMLFq8igwXWMMOe8pkaUcmIFw2iakNAiXt1Ag9FYzomJQADemLiGe6p
b6N9bEM5+uq4dQq84azoxwlta+d1DQGcSx80WCwWjqrS1znmXvK/hz+S6sM3TBwQ
7gICm8Z4lN7S6JgsFxM8mTmBm6N6q/2u/VKaChH+un5sW/ZtDPVJvD7eG5QzjaXB
iPHU797mPMlgOyo8nmgmQD5YoRtEKAO06d2dibBtHfnGgoN0y4ZGV5m7jG51+SqS
lHEtATkNMl9qZEnwd+Db99Nj++WC/Bhejb13wUq5qzCjsSBa8XgWoUZo5t4CrCBZ
tRDJmu7g7bAjKE43n9z/Jg5gBOvlDiYGm3yQ7QVgO8t7IY+ag7quC/2OzJV38+pt
0uQqcVLQvXkEjbiKxD1YKlWdSlf7agk15EFKdZjm5kOOY2Ml8DaM1/8m9W6qpk2X
myfp0BnD9faUiaZgJ8n1Ft3vZkyjnVLUkEW+jZqR3lk+s7Zx4vVnMcTjuQH+cvh/
PXEJqHpC9hh8Pur/z8JH5HMVVyq1+HTe2USGH0LI8UJIXCJKywoU+hKovwGR9v5T
+eFG+A8+dSQmkEQKQc21CwQGeXXFSUntznPqEAXKY49mPHRYI7HzrHqrezxodgxq
jDyhiVtWargtwnQ2RQlL8kHam1q1vL8QbdP7HU2tl4POWpNg8qKQA7yCMwlUBWn/
prWtPlVuAZ9Z+BXd5vTz2tUxYFPRVDdnsK4lxg4OnINdiyCTZHyN19IYM0Hv0gyE
e/qtsu9SwPZgdaohyMwk2v7+FqXBy/L9ZkiLnbYFI15bTfGO3JTf619SDEWdzKz2
cBzi5yI4VdGHpQVhneFvOf4vRs6xkjSojz2rsb58bj24C+fTYzc37y3OXhW7NrIP
4M1B/vPw/6tnWkRhfqLOce7hCJZk+ojnweZjpc+/yfTF1JHW4Aa+yCu/DCQ0sH3j
gdoIFwu7AbLNsZYDgoYJohy2STU49lh3ZEHYctpvvGuWpq6h1eT4HKpGBVIkcBcX
ZW/tHtvuB6YvcQFxq7vP7oHlenNESCDRS6ixWcr4B+qL5MeyZOlNK9UAnPopVKpf
V3oM1QmFAhhz8d5nyznOgKx2BYO2PyoZGDXbDjE2X0/I5Sxn0GgihuC/YPwspKj1
5dCZSiAS21HbUszZQKVI9Kd4qCyYAKMM2zLe+LeMIHRuqoSEd1bn+ZE0XR3GeWGz
yHovV1JG3QXOz0WkrrOSmmpDAfFKllEtj3mGG23kFc09mbhVV3jdBKs11YLBK6mh
Uj2lZCZ9qs+sG5Jz8uv+2J9EnNzL1WtaI7ukBQVzr6+nulTyGoEhzjk+lcVFYrhr
yFOnOAPJCyUzPTj3nrFHpDhkJG4wl0wMIt6VdhU9b4IoKdXWBqDx+0pUDOoPS1JO
7T1wsGShz3EhaVuYpuB7Re0Ye2KqyCMGASjYMAa8kncDLc8ym/B55+nTaLFD1fEH
Rg4m5At/ZTs2q+bdWK6/PljHQm/v4clZYhyDBaKaqxjOxxqSQE9YDygWkgAzRcpW
epEBGmBHGqmzt3/WpesVM5ntviZfO6AXM1F+CilHuLqHE16q3ymmARt5GX0DNUS0
StPgBxrUhajsW8R1goBHj1LtLUE6gm4dPyjQQiKxGd8B+xFkp45M3ZkxlnR818Nr
QLoYWHwf0cdjKeGfu9K5dEeG2TNd3AoIcjHi7zpeTnaNoz2fm9to3lrAtLFV+v4q
7WjRzQY94odr+1p5SgCsUSNM9NmiMJ+Y8D/MqubyTn2qwsRYt0Rn0lj+pz9H8aUt
RA1VqUFyoS4G6jbwcT10DRNLdS7IB4pXEc/g8sCIP04gJVGvLUwWP236/jbN9NWS
NnY1SUotrgklfbVvNkIIDTmU9zDcf9atgMm14EqcCS+tQhtbB+QvkoYmvPoXO5aY
K2utQPkGKQH8YnOSAtf2LlLz4CjcJWFKU650S1nexqEbe26z9AY6Y4aWs/ONxPwX
hVf0XtoCy3avW/tze6DB7AH9gkS42aCmy+f1U67CoI3FWRuW38pOpprEWd3Sdabt
bKzxRI7U9vz0SUDy9h3//7GkvqxJzhQv4wzl3UYieFx1qCUzqUrw6FqbpKtr9e+m
j6FhsEMGTMZMxo081Z1ioDc6mFoFExGSzIHvvW7PUjgc3SwWtFOD3zK68oigGa9V
75hG9wrH57/3XdxvqsznaEY4YNi+KVZGj8eGEycVWYc8k1MWg+6K276106HJvjqz
HS183p+gQ1wF3E762QiwZhPUOJAo2+jxwsm+3BFKwpymHA2CyP3iduhWYWmosAp+
eXwRlyvziiQZKWjhtmUf0tNQyOrqmYfSV1jTiWxu26TyHsNh4TVgjcTLMLE+5g7t
uduHGHu/YfScax0FYEx2FB25VILRUU9kA824TjvguGi4LQCYOXz2piFVMjp7fZkI
yBg9t04zuQKb9QppdWEHhDknjaiEaJ8aU1WnVPfT5t0U1niutzrRHNdEONFlMuez
8uQjQEtYi079PlKwJome95Yf43f+XVZ5aQ5MRFu9CiWY7XPV7zpgahlgpZKQXbbx
wp8/TWYSO9bbBBEZO9xPhGZZGf8+Ynl71q2Zr3TWuxmtqB8qFTjgj+FOO/ZAOzrB
+sY6+wdOjra/9uut9lQMubnejnt1RK2KPhx5SkpJjy19RrABIPfchZY3Js35tn9I
9YMKvZWBIpvyJnzYkdaXgCB2p4/ae0PvM1hmZcn1xpie8TgRW+rF59mashoCuBme
CYwWlUz/eBkl9Iughu3KoxLExgPvTCr7RRUnOYHvOADs6Q4UYO6qrQJWJaUs44EX
AZUQxolL5DRswqSWGKpevn5grdcHaj0fCnhqspwPpx951xOk4hRElO02T2awkw3z
O/F1RGM0DVvCY5DtaJgek3RdtRIyWpjOa+Z7TkBaMLTfvmCsgJ3BufD2RBazLD34
OsPHI/wCeIJkrO4K52QJl4fiJxnfmfTLAwsgNTJBK+gH/nOmtuE5BAKr+OXbJe4i
cZt0x1ti/dmxweIG/cEPCWjg1bt8MOLUg8PStzMPvTMIBF3jVc819zy4h2ZHB+wR
98q0azNmJxyf4zWyy/BIsQd3OjQG/NE6rR7ZkZszCk79OinikPKDoc2xqGXVQQ5D
63peLVacrfpY9Q/WEiG2c9nNpjpWRHy8bYGN58cVYaW2O17trLRS2/XWaV9Ob9Vv
wFXIQn5CLq7Hmh0CGQlcyicPaUAi9EbmUQq4yhiYJIO+jiuH6trwAHP4C/ZCIECx
1xcJr/nUEka+Bk7011fVyS7Rp2szQPv2onh5fFCY2+U6mAAlIr1r27V0/WcQso21
ZB0NXz/xd0LE5ce3AwjB8kphC8xg9nu2IBbPaoAEyXAZkk0O5yZr//enM0JGcNby
8En/wK4G+GrHsTLS0fTTX31bL7/zlkRn4qVQqvYqXu/RxfV6s6poUsOAyX4pP8TW
Jupr5rLXj7mudjnhWc61Avg9w3AgPDd0MwgKiJhiMP8uuK4RLdhuPl7euBc86CJP
/A5VGEUO0K1VTAMLgGDsaABbzfAwGWxZKOXeCump0FcA25JPB2PZ9J4nvIL+Zyrn
G7WyGFrZLZeoSJKOGy3RfGIxm1U+omSZpal3R4IKuTNtOgEmWipcC4nF/RUq322n
pthLV0nRQtdjtrmruuBSzSzI9dPkVowF96pDiFWomh4ZfG1BOltsi9mH7jE5hiGE
RUUq0b2vtL1SIO7hZL1OC4BBVGmPu8Cl9XLPJ6+/gKW6duF8VEicbqGpjwRBIr7M
4lmzQgrfkZXx1RsCiqa4eNvi3Y/Qih5pymHkeh7MAH1tD5ij9MpD5dlVjBQ4EfpP
xjGMNGkCcc0QpvgbAq1p4G94glTn8+/T9BAguyITrEOxHMptdTfybTazyIeomosn
yWFM/8bkYxgstXjVvw8WAXz5vdx5jkHn4NxIrXgvnRB9qPMSRboDAphkcsWPTfHb
hFhLF2Vip2xhxdHEoj8A3hc5o2W8T9zCpylJmt5zU0EXcZw+Z0ZbZCMsbGmJwAIJ
cgPEmpy03OcsdVVKHKHQXHE5ReAJk/1KRCbeu27jOmgCvC2wCK7UmOkKzc7xxIxi
hzhJmUsQ0pasRzxfxVdIgj0soW3ccqL5d5ztuR8F0y+WR3jUTVdTYOd2SQyyDQ5P
cojbVvlZ3Mepkx3vKyvj0b5UUaAWWOagaoXRfcTOQDi3ZQ/fi8ggPnMxRJ2aOZvu
iXw6kIpL8uSPn7UMR/T230xikYhYXI+g2HYkGaEaUwPrhTXmxvYCfOYse3RlV79a
fZcKO+QjQPNCjc3N6qvlWl4Dti88BBR02GHS3He4Bko+PeB0Rx4CT1yVd7z77L9J
N6ZPgDIsq4/y0yMY7YLJh0qwQvxZ0j+p8emQbNfdVfHJnsxFecEqLrSXk4usQTz2
E+Uvw4HHalNbOrbruo6LzLM+0bEuIJK1x7k7eKkgBaUFu7hrEdPet8qR4T/csXxW
EKWyhhClgI6o8KRX68rd+F2V9DzwGJdn8ewRso2nJX2xNgtmGi24cm90+KsIKRJE
BsA9fpIfzeCWvFvaREtaEJrHgh7Z7Hu3bcp8qQN/tlNHJNRzl2oU9B3VF47x+lyf
/nf2fjnixZ6mZYQPBv9lhySEsY8HOR/clbkOkMgMPFX/+DqcHw4Bwy23NgRgMSy4
XbPk4KVFzp+F+9DVPSVaUg3ujmnWIHS2Aq1qo/nVTL1lfnEV9mRq5oNG/rx6T/rA
eDCbKF3zbRcHlqtoeM+L2UyUNprARQgueCThssSwv7gxgNVuZmBjJ+DvVyqBIhN9
zn3hgzTFvRHuwmp7wTmYr/sZxaM2lc0pgR9xuHr+KXeuFs3pUyhfBXDizV39b14N
ZvrrKGatlaCUIGl8pheK2q8NMqqIxRhWwLsFHWibG0ltSzFXI3GVT0Q7cwnI7BOO
cpZ2Hqlp1HZztxRLK3WTZTlDCvdgBFwXsDlsZQC3uUGUz99DvhHhUkxD175vOoqY
hvJPZkwWgJTquqN1Qx3heAyNBVvsZSWHAcc4nxc5OWlhPFHekNwIuOkt6iNoc21v
VUip+QgHmKivgcM+9yXGPHC25W5o0ex4SsmFNzGuyiniKLc0Ll0GVFYQmPzdeFOC
BYrURuVtT8CYlMgNI32xCfSqmO+4k0FM0qnhhEl+sPhJ5QzZtHJki37sCK85zvW9
lhXJ1UrrrXQX2nAczGvRtg==
`protect end_protected
