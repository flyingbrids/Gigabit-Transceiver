`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FtnszLTM6ywe05YlxRCPzRNeKclota+wn/WiPoyyf7t/E4fbwhHTtWBXK2gsaEBA
xCimnWZpAgeXEoPYBw7PXlgEIGjUeLnovS2cVyysSXpUiDH2dLz6YSiU8p0leKuz
eyfi1ihQWms+hg6IJusXCkWm5ZkJ7LN9l7OqGtEcL9Df19u0lcFeMEaTfYfsYPZr
SjbwYrvukWqsDqyHkwipkwQJ92mSDojXsYl7sDwIxYs0ljzzdE2X1hzUt+kuQpOI
4RQzOeFlMYI/ee4ET2aNgLZqzuwweMQGKRdTD1x873iRh0UCPWq7L9hapz4tOF4d
XpTj9YhQXoy6qllJUNEL1g==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
OE63U77IWSAIH12sPqcCr0YCPD/l5PgUjPHxrECSoKcjPRgUVQEUXi9rpXmfAOuX
/Pooj/ZJ0Mdme3ZJGeceM61bfC+FoGobjcHl1uDVcz8V1LvkFeIShDFGQVRHTyFm
QqqhmB/aGo9GqH9uiB0UWkgODtLEoH0vaYpCf86KIoU=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15168 )
`protect data_block
RblIYOo/t06ZkIpztpguMuT/ZTKzVJ8LZqor+xeC+inr1574KL4No50zUqCaemAg
fKPXDX016gZOsxudzgkgXOyQ3Pv6/WXzp4FNrU/fgzN7vkXosB1aOyY5Ym4M8FoC
tzTG06SnOr/zO2BCh3FU/KhQQVLjOL+ex4XT9+Mv+W711bWRFZh3FqE02laOA7OJ
vsa2vgReKBZ+ECvUbt27rhqj7SCJIfdIgRRbUe42wsRI8rGtunF6Nbl1b2YprvSs
LMk/DJfUKeQ3p13ANON3opf4MnKU3xi/DczmSgOAAGHJSgYnrtI41nB04alZNl7+
jQFhND24NQafikGOP4RmGNnZKOcvQKxCZclRdug3f4Xt4CdW3M/UsHTwUyRD6K91
nOVhmAmtrtRsZaej+SfgfLVWGEwf0LNPk56UFwB1lUJ84vlEietyj5DnBea5l0hd
nO3ZlaGUX6bqdoPSsr6ug0Gd5Si3bmKkDtd4of1qNBJMATOgsGsIU8ZlFxtVERFl
6s9peoHRQnwnSK0nvLq1G1qB5ch3LExNT/TkTshe651Re6QU1AB9vUniI6MTpIBQ
QQMh/oA5gWbyGmmmaePiZ6LDGcR0Jj7N1WzbtxfanD6A9sZXZWRaHHmri2BRQzNu
R7m/tfhHBjWCShgSlmdL6wBwA3XKXcNS3uUBsM0badEg1qZqGuGm1ZlC8vJlVyJm
xUBWc30qPBSLStWsTJ23wc9B+FA85No80ISCh51/ztbULtQMSWgoLBAtpT8uwLWm
rteVbT0mmw2OakuSanjPVPiCMS4E5uIzz+pLTXJneRd9uPL1Zga6hVEH323mufBZ
Nt617n7AxWwP+EOAke9JJg1ZXeLZTkDSIk0nH6/TKJ8sj304tkGPB6jCzbVkjSLW
Takdc+vlwRS9XPhcYluFB4aBDfWy4NsjZigV6eZc0m4TYquaQamzOCJ8gnZOx4e1
I2mwac3A7xqy1Q8Kp0jJTR6Q+oU4RyUGLw6UyLaLl3OBHAspHz0qZZz8JTxgvmKf
BCXR33Q/zfoUuVaGePJlycLSyiKJMQUYC2YGhWWuVrSxhsxBMSHpQdgMQHYBz85z
YeuetCo8zxm2I+16jXiL2fpV6NrqX1YM9HdLa3HJ/4B26hLqlpibIVLNA+vmTX3e
ovuAm2OphLms9LCAcJb0S9AhIPThQaxjziSzhVXsAQ3bGCrKYhoJnpXa5zno0pK/
QlrKtKIv1ZntVCDTe4aaaZvL2yqRYMPSkAXq/PiQcg60S8oG/SbfVGlP1e7mgxsL
d/YKAevmHnpI/y5O1p6pXOPR2iSH3F72paWpfZsJ4SEHsLs9pxFGpAQh6xnuZtLX
luJN5JyMiRjatzlmGbI4q0P6IGMNbMs9w8uU5uqfz1cLOX1lZGCNyRbSBL0QCuoj
2khF2Bs0v6nvdQGO1qvrLSIvMA0iIQe1S5RxDYcAE5gDFIOYwZDxAXQGoGOvViuB
G5NKAB/t2g899RyMH9b02fZvAYAKFBob7FkxOpqycL/qMgXehG/ovUrGMV2lRg0e
vKAyqBRUw+PlUcav3e+se10TOjd1kL4V1C5tFY+/TNeY+gnUlouY2OiVWOHym0bq
tZE+Aud6XYM8D2eN1nXA7tw0IdTvSQUR5xok22qgSfLhJ8M+2Tm9Mro/0iXWZBST
WqJYdTp2WMUX+LsW+ii8AXi0vB8d0Oni8JiHGZSTO67xPgqX7sxTgTKxZTfn/xcZ
Cvivc9KIZypghHTkCdSYiSKWoZMZvRZ1PdY7QvjcgL1xaG4GuvlebsCJKL7fayeG
T/cx6e9ACLINM+iRi7Ru6M31vLcvmH/mi2smqvEICFdmRTSYKyO2fO860nIKnwBv
2MZx1lpuE+Xv8i6RWtUf60SmlLc4q87yYf9+hmUfDo25vRQLDBFXG/8Dcr3MJcpG
T+SdZBhA9d2Wr5JVmUO7NWzjRUtz+kSwJpC5FdG5eJLGKH6tqjQxz6Fg610cVL2d
SwBHHMk0sqMNr56pag4dF1xG4v92HAstqFDcoYd1E8KxV1luDuHWM5jCTL/j3b7w
ZlS/sQMjHuBLsQEUk7jCoj/3VXAaqHvp1SkKQryBuqRh9j8W2Bd0sxn9307QQg4f
V+EHrSHsK2tyOkGaoq9rjLhl5fE2DxPDDrC1BwKvMiI55aUbLwjE2P9ha8HpPz79
GCL5+HX7u3shqYuceZOfCCU2kFwfZVFt2RlnIQZ85q76I+R/hke/OQ8qoxfahSTC
4zeMGibj7N7o3h4PBZlVgZ4EeOvZox7AkrnVdz0HgWUtjx59/yod40PB73w+hR5u
DuAIljVf2xCjKxBVT3ENbqpotvKMqM4msyI2Sl2MNTaG8nCazCBVCsDQitUCZ7Tn
KsdoGIx2DMiLeib68nWBvhhpo2sozYnzSMhfG+3lfP/458JsakaKqVBBAeHjRBla
CK0eizd4qxiutPZ2qwYgOoFLx3arZ25aYGoYTeR/xAu4rAyMVfHIZ98H/w6Lq+/N
CQe8VWnm3vBBM0AVxebDcMNQ3aO0Ebg7er/cxTrX5nCAjdXEMYov18RHV0sdbfSK
Wa+eeaAYmrh3+l9VgqGte+7VPgEZmMAQAP+HWsW4uFHVb6Wxe/UxkrAtYgiYKUZP
T5/DLk1mZTCCVrfV9M9R01D/7qMJjgABCvrx2nUyyfrAM5OnB/HDwd50zvY0m7xP
u0KF4vYwNct20FB4Wjsn0C0UwQMeTxhAnwPFfnq0dIEdJf/yHW2f1RG/CZM9JMHm
LLxEUD1LSNQbb9O7N+JD2f+19Icn/+DpNfqHViiWLt1V3vN8Cf2EbyBbHkkKrUG/
OTSUC1kMbICtHIRoG1frBoxAp+Te8lzkBDrAC4k5foZnC8YDmOzYIwtWEucXtPAU
Ob0D34MXG5hTXdXg3ufN0biWTHbCi/BsrfbbSeBKjM1uTHGgOr5+6VF5MtjwAqIq
KjRQVN7MtKWmnacQ6123oT9AWF5INfVxt6izhIcNTgEi0JFt4LYudOl0vhWhprTG
b4c96tK3sckwjz2vqTlJJipqfRzwrQFkUeGI/s4HADgfA+GMLpFVGvkWfrDTMye2
XPQCRMQD6w9UW88xkAddTjt4WPItv5GZvJToU0v9HbZJa93Cg49gilwkyHgWCwoT
BNEsVxWEkW43ZTJpMqn1d3clLpKZFeyezpaZI70LoHdfVaVmsjDCEFK2r55ZZqP/
8RkSUWcUYrcI/dWtLH1UE6w4/oNErG0Mg5ksw+3Z9SATaj73TeAG59AWd54p3v/Z
SOSw5g1vkR+toMowiwJtO9D+JNJqBh+MfSNtBN+ezrPLWU1GW3X0rcsJbYBCBotd
9HGdDx6WHsyjpJG5ODyqVIYOYPO8Oa6DtxYMD5TK3VJH0IP8OZ7tDsufDTB1FKZr
f5uxGJWaSTVe/xwWWSdR9P3Y3pEWg3Rgb/wdI3Fe7qAvs+rIt9tnsCs3TFZv9ASQ
Fm4n8NMx4jK5p4to5DQOimmL54uAk6jZq2qQIzQFiU4glalAtgMzPKCRJolfNsBL
q4onJhS2+9bEzJVJ8CFmjCkINAPUFM9/67qK1eJl0C8XS5zuG8n3//zgz+aK/3LE
XYSeBt4lrBhYkvvZzVviNhVKPV7t3ckhfkgebkkk+eP29elTMI3/P17DkmZz0CJw
QnpvANw1JfUesKkxdu3MqHP9S0m+rRUgWFfH2wHjLtQPSFD49gLWxrBGbXsRYabC
VvI8MIcYrLJa+4M2GQSnfmSrRWoVHGCDlxH2OYudjpR7oIyWumTL4oWV8R5dr+C+
Ao1yofDa5Tgj98r9K2YM3vZAk/oZjdOSFZBTSW2ANBoCAVfqLU16YbGfAhJF3Zqm
bSyx/+PVsM2zJIqA55IjdrpMeHPYs7I52NcjnHwMyKd7OVJWEXsumTIgksuXEfx3
NgtnlKG4+d17A4Fgwh1EnlGMzhJYh0K5E+r/iQX2LmdcBJHYyBSSyHnLIqFZQfup
pkaGxT3qBbTE0kln5E68tQu8ntTWB0ai/xVFWQad6cc9waKLweW0XxmkVEieG7ZJ
L31Pjs9xhyiykKoLoeYPPqSxauGgES2xjUosEeURb7+oqzk53djsCesk+pZ34/iE
chl6+pFO0r/TsFRfX45ku/608H85hDOPWxS5KpV+kksB8/ztQAl55wwnykl/6zzA
gEWW7kC1niTuXsJcpoPdV4YddnALxA3m9YabQsMtpJo8r5NvLKKep/PsxwQTLEdj
+FDbEYS/jljMtGsYV8dS2KZbZfiHGMj2BE4A67/4NdAxZrVVOEMtjzCu34RN74wB
hPT8CJMo+Fp+BvIxXZHoTYbcD9TIR8dGkKm9r4+aHwDZ92TNAwRl7aPUeRMDzPZl
m4gX7YwDIwA+ZQvIbZ3Gj4+b+joLV0B/HsGAxDC47TRDlGHAFuEe98C2uQFeP8xr
XZNJsHWHr9Zjm9EqXaeUgWQcK0hWJKMfCpYXzOrDAGHq0b9Lk1jLeezBho5dYngW
4MlsaoePaCnty04xslF5iNMiT7c3jkPlXOrIpAEHSutLEnKlYtaTD2SW1NZ7W2pi
zJQc4aeV4Bn8rYqf93pf5wBO/kYWWABqpbMZT7/2JzwCxf9dIwrtuIGqmE5eJEP6
9jJ5/gvSXLvyq89m21dYDm/prVaUvHk2uRXZLJqfftElOnWnBSj3fgDBq71Nl4/T
T94XOp9O4k9Uk8lf30n7fZTLIjq1SZWhiyJEWZ2+K+bMn27NrcAqOJt6hY4ME3Rc
m8rVlPbi5q2KYR6e5lFlEYJ2AUFudPYeBPQttKJ5bMCpFS8JKzZNFSrc8iL/vYxz
+cRJqGJsOOc8ro6UvAQ0QHnot0SufVcssS0T2KmIsARSkRpeh4lGUch/n70jWqNJ
uf6TyIo03ycEN1RvtUAvn/HtyE8/MBT35gsDfwJ3sDkvoBoQGunsxTbs7aECFNPz
yI2Fi1VEs6yt43DxIK0aA0c3B1bx6DVzKQ1Pp1c2PH2hWMV/xBne0nLQDK1Ao3Wp
C7TH/wPLagbqK9qohExUU+Ejatm+n9OjwHOkrQwHnShz/FMw+dn97d5nXFOPyFnf
sKxLu6+Tl48Eef9C0PI8mQB01+QZQN0u99+Z8wUOQarQWiVtsB0u5aABIfjLwDAD
71UfcnppB+OQcrH74GOLM2VCI5iyVYAboi6G5tEMNw0B9lB6Mt2hItwVSuEk04V8
k9E3l9/O4+I6fsHn1ckWVFrCaU98VpmjsJwRtHXvrwjN0xmd1LFylgv03P6YC4Di
w81L0UtCLqxNjP69oJQ3jQYCH8zhgjdbF77eDVP3cBdDS6FfgHWOauSPhooSBxF3
cqoGgP1dAnoaMsniWrEeR+IzhJInwlvfh+zDzfSGl5e4qJdEEaj3OyzF9ljrBJOE
tcg2RLdo+OoQ9Z6e45KBG89GuxeRhGFv68aYMftz2b6vRVn4LM/6/BdYkKemRNfR
KqDvvhBUwzFdCefDiNOuVQiU4yNqyUXau8WQyeQFaTUKpQOedCyL71eHPPIj+/Ik
Xb8n6goXksZydQwilB5e1HQcYY6hXNjUy+MWcZhW/PMzeCzY+wSqZcE3EwL8dRnI
Ag5d7DsgwvVbODbSVrQVrO+DdoArTnPrlTqZ6yPGchiMlRJVB2FT7fM9eiWR8GdK
Um4hp3uCl9dKJJbSQTVChYueT81+XXBFNh/ZDl4pHbQmOF4qRoLtDq9mK+XvvIIV
2Qm9Uwf5YaW73U6cGtdqp1FZvBnkxaDw4+D1I078+vlYipVFNG47Ol9LCixF1ayp
AU7E+zAFWDXerIyi0CpG4sNhLf65jaWwdKYqW2yINOesOBXTsoKzsWKY1FMz+wHM
9z+6zpD73yEi0dQIj/UnrsfGRcooMJ8LlcLvIH5b7aG5RlRua12b86MZZvYusP8Y
oukoSKQNcRoGdPFK8aa5qP0mDNhiEQu4rSv95Sp9qyMKiF1v9TZdthMBF5mcCneU
gHb0uzwBW0WVxdC6fOgNVaBJDewHjPxJ4om0MUOMr8x1ktnKoU4esV5BnqNQGZJm
xjb5UJDz0jCTHjnSMGletF14nRHWGyG2hDHgZvUd43I1ovaK4vg3bcmnMjpgVS0J
StYsZ1yVoGIlBJ5PrLhQZOk1KcAlVC3hlCxm2KwvpZ8j15NIPqDCEOUsEvLTqo7F
JrhLZ7B+/hT7x307KzGzqaB9oMCDcT5cykqZKNgvh+u+TBfA3ZiQ+W2RJANXZj8c
67YFktpD5+QPOEm5pOb0oBT9Rjd1vIdmeVxCqJyPtG2JPXoCrGP/AHxHLT209tJq
q/vxfvlEVD8HcAsCisJBHBsHXm2CtDWWs+25UTJeK2I/MpNDVQdyUqZuJhHgrJzz
IE0gAmHwd246Ywh9NH+Po/s9mhfIgZqfhakh5QHUgLZauXv67xZeDbGSd/9vNjzq
9Pj5d9c+1P2VFSUVaBTcn5crGgz77aqq+/XmAEJjauDfR0NIbUF6WRtjB9PTo4gW
uV0yhYuqshVF/PR+I5UH848ucpVn9NfB2RjvtSymc8xeKQYo+EZQS9oA3KfZxmq5
MJwX8XjRuBTE0DemY8RWvKkq87VrL4us6EoO2ktBRP1YTqJSEXZZFlvY/IV7j+4Z
R+Sjy8VYZd5+YsT1wtrPaRiuNnj63BJ+7NUq5hNnLNqn0Ux0IBSAR9EgCpku7RHv
mZpwyYzrSwiZ+OxuF0cddhc4IU5iRmFn70H/nXucLxYKDoOuS79RlzN1aM8Ock0Z
bfCc5YBBBhcknS0j6+B19ufqC6IzZxtCiyRVPXVWf3eHi75jZJGEmPaef16UMS7W
LCDIljeXva47sZgYdBa+QPyOCrZb5U9YEuUflrhxH4Kk8Bcs6S0iBBy8iE6Hg2XT
O02iTJM0qnHSu7WOFpQANnwHG9xcveiQ0hf9bXuHQyKxXV5RX2d55Ji9crc2cNih
PuVNjqeeKbr0qA+9urSYrOZDUA2tPbrg/pRBELIfUYq+7z3/V/O/TC91a9wHW/pw
CfUfolU18KDpUdzTjuRSt6Vrw8mLy6i+ITpWvnVaR2sBXwxfNezmH51xEpUW3X7O
tHzkEe9b55OjVwtMRmRdrwCMbV6FjGehWuCpbRlQpqHFdz3qSN4jBrp1aFUNfVCN
pYdnKOUjfa28NzyIZhGYNOEKEjUV7Is859qD+UmE41oglPJ1LZiGW9Ct4nDYW4Du
IzyumWxnAbtQ7e0SgDwjkx6ZSgj9ddOw+7AXg+CxIzgPV80yhM4e/y6oyPTwlS3f
w3P7oGu2FoTQVX+76nea2xl6uY9XBHNl3AcPTnFDUqzDqSXgaBS2gQ8QZnZjYYqs
hoUI4DGoD4mF1ixaGJbg4KKhEZnYownN7QCD5u8pNF0qP8dKxznZ2eX0q3DBh/y3
0GrOA9QpwtxRLJOAqElSQgtZ57YD0bJq6X97/KKQdgR6xAhGj903q2LxYTujLR0k
0Jgxo0FhyHWtp65KWDARkOds8VlbG+9zanE6MMAM1VFTztNKktR+k6pT9a9I0k74
3unpQFGW4ByZmw7KmFgafUKIItnz5XW0CprwpM0IHSbUQ0O0GNH/1zKLSko3psOa
8zxFK4U8qM9FYsU0a9MmB64LgVMjKtcOdjpvtBEfp5h2SMHUJ2vDpiboYxm7O2yk
3p5XslhMo2A2NYXxxYes+E3+fZ0yDxSHJWKrmI8gRS9DHYSJKZ+p+uLNYELkMOod
b2qJEblQEL7S3eRl+JWgbEUBCTMNzYcnusV7mC8BAbVQIfD6HLiO31CqbNVTgEzE
18iRIuQGBT4I/rZMm2lItLtbS02aeKNZHli0+0Jjv+33u4w0c1uBPKlZcgcTT3ns
mhEHayECptjS4EBCS/Ob1ogcuKkgdaKz4SKkSJSLS9nSWfIjohndxcwXTw4mNMWo
vPjgfpWW9H/1TmwOFB/dkKS0Ml53avutq+JEG4YufW4Z82BaeowihPMJUeLpy8Qo
tJ3+MSzzusjNsKlgCwkpV0GIOgyphr4t3QwtBe6fn/O8NykUAap1OpbuNYiY0T83
K1f4HUa7CEjoqQh8qmnB8mGLQCC1hYZAc2HajleKEZezuWCd1Ko+8VygC11BznIA
Q9Pp+k9RemUb0GsR9CQep0j+AQuwzQCPhyCmbLOYXwzL7OSpwGy/EKtR55TzFb4N
cQFQzOwL8XErUDUjqAUVJi+rn2gRnyn60Z8Rdt3Dzjp50DcCXbKSGXFsC1HZ3nyF
ixhOlgjRo09qyJbTUHMFva/TYFXR29izmrONa1pxrWNHRj4VfWLA4pvCD+nXy0fa
o8Ox9rSrqT0nAdEwu1p3kj+DoTq/9uGoxnfc+2wR+TIWbYfJ3jDO8+nSrx1/lI1Q
rxxtmogXJ7CY5BYOkwSmfblAIbo/vC/X4zU9DjS3TWxSu0bwrgG9aq9kz9z8WHNa
GubN9+z3DoDtrBRa2adcaAKzjJhU8cFWkVubL4SscCeHkcayJeh0B9W+FLhJ6U9I
U5tLCwJ540PrUJAY4tPfPBDttU26tu8AQs2xjgzEfuwadL7AS2jy+ES9/1M9ODG/
UwEnTFZV9xmLc9YOX7TazGgUnoWrOtf2cW29hlYST93LuHP8GH0PsOPD7WI98mdk
YEjyADpcN7CZ4oGIrAlb8WRis1QOsqKgFsunDvH2JvMhYKjNLRyrCTqKfIgr1eRz
L1SPFMnCfjHZ0T10CvC4Y8Smfmo04oC3WZtpMu+6u4ps9MBbQri2T8GCnMAvLnvs
dY59hptIgfLg//HnzU3J9Jyni4VfgOtD89t4uc/hVAmkqq8T8PLoDtEfs9q+olYo
8whG789vKykTY/w43yBGimMH/4h7MOrBFb9oTn4UYqS+BCbRYciY3cR17KKvTlOa
THu+tGTPbvWYzLOMBeguaLZDpI3oczTDhzx4j4lp/7pfEO78c+1+SVWVIPnLe9yV
v2xwHVqnK0u013NP5nqyJDfE0YOGYAGptPv1xVF1A/6L0/2DOlEA2bmNYTqt4H6G
rGcnRFuNPI+Vt17WcBwn/VxT2TjvM1B7SV3+7SKEwTCvfoppuFGua67KL6yfeFZL
7dEuoTRCEVRxIOpDCEH+xOcvmxDbfKn/jda0Bglq1c5a6RKDYV2/oLNPGWhfmuL0
G1hHX7nWja+s6yuJu7fGb+ch1pbJ/HJjhO0uuId6jq3cLW0WOPXxAXeNpr+bv6u9
wPMA1tfeGRHoXmhHf251x56JC8BA/8k2LyGDU9pogmYTY5zO8oE2rd6aAtB4QREE
94xIUW9o7LkScHKzcgPnlUr2gZ8PuQEic4/tqmLENheLGinP0teJIvmWTzPRLYhx
7ahEoCXkzbeJpVIwRYFz3WVaYHQhMtnK4m7Zgk+mdfV3kwsX73xXOqDsttA8WuKE
x/jl0wU4jwz4oRrgp8cji9moAJzqLqtkInqsnKGIumJR8J4wUcPLvmx+ClXuLTIv
3hkqezJd8Vtc8FQFJ0ykxj66FOlSD1TJWA4irG1Zq+tW6Px8G36TtI6cWHiQVv4/
sSJV6K5XfkrAQTBmq/DMbPq6CGlLswE2IeLgai64QYioHOMf6bkW48PUtyBYFkcX
j8W6GfNKaG/NTcDItaYtppzqoQgs6yWSmLvMXbhvWRiOwbJtOMcfmjz0KoKuMGHL
/Trouo09O7b69AZeUT9kvwT6AaWWLYCYV46oYwkOAIOej7ZnYKS374rYYWxQXuy+
cbArPrJHk8B9LhIOQLe8V6xrxcC/kPHfad2m7Bfb3/j2Uz2WOlBv7AYFVQH8W9s/
3DMA2FzszLhJv/8LIj2staimVnDPzDfh2GDMaPnSp8cASeFZ/1o0AX9E2O4CCL0r
IDDsbs9QHxEdBYudfwHjlHIzLK6dIzBXgksiCoIr0pDr/ISHgm8SUiOysxQTUvg3
teCqa76Tb9odjUXSDCnUa6KTwt/PJgRc78zG3SSnCqkd1a8o1nnImTvs71et5yhl
WCD0ILrMAl7V+XCHhQruj+oo6XmC7ylFleXl4AvW+1+xP9AXq8RyJdfEgvuGo7Hz
C60/lrTUirCwahiW7cJ2VTLPOh7V99QxUsVHPZj/yjH8KMdFejz+XnPAwFEO/lZQ
bqRTiDeMgCUpBOoeRvtXMXOzYOnc9qlfc3b8G2WeYq0vh3pX1tWaHWQrtlw0Zzrp
OPQiA6+Z2m9DsHi4FUOZu5F7LlG3WC1ZnvnxySkuvmbmYTUi8rKRtGj67SS8WqLj
2+927EBnpStU4LrHJ3cGDma9hGkrRw7nkyklcd1tOKm6gDDDmQ/KB+n7NtSWezAw
eYUS0wRE57M/fjPy7W4DVNu8f1HVla7KDcFS+SXkMiUzHfCLWay0tXuBYKTi5VrK
TTWfv45mTimqgbkiHLR6eUbDzrxR+Ke2chb2ld3vwva5jg79HWFXQqXfdj86LVkq
7V9qTacuU+cRs1omMojoilhBhshjlScDuAxoFBj2tN6M1oI3NlcivKEgdWd6hLQG
68of0Vj5uiR38WFmy3tverHgiVG3gsZ6V6rdBNJ9RKje88HJ3ZG7g1iFfDCIeN0k
JO4bAbKaTffNj0sH2fRoV7UFi06E7VPy1AVYKMvTTJDGVWWmTN1WN6QIYg+9/8OM
KDrOnNB0nalh4Jq/Eq5xFsQ76aLSNQh3kjo9KW4dJuT7McedBj4MwoxO8zuO+5gS
gWZmEjSdI2Z/FJw1N7gTPj8gR7Nwtv2GPecqr9wjszZYeIT/OBBl8aoEg1N/6F4k
s9Lc5ZGI6Ie8UTmds0mCXK8HD/7okTzB2Mq9NLkpPw0h/gabM8HXktFpgB/M5VZ8
wNy9BcCAPAjS0S5FvYSTQas+SwfGwFI5cgnr6lQaStwxDiVFnj9bQLW/ZQyJoecc
vnXcUVAW5ofpdH6ppsvGtht8EeGYCystsMfLjTzI7uznH2JgwMXlCOgd9KZEAND6
jxxZLHv0Uae2T3jDMt2O4HDpO3RwX1w6TqVPw54VV3trxsGrLvrE+X9kkkxQb1/0
N47MTCUuRGdmWuH5nby7J93HTjfc4lryPD7zh3icwzLzwD7r7gZo8afyA5VhI+je
nn0pXzlM/WfvB/tm4Zqcod676Ey6gLzNpJodoYkbOVZmBAd3IgqTclhnMRAyp9NM
5zLKhcDRUfq1yV6VsNVAXLTS6ZYr4+S4pXMTBrOOBo+wjZ7HE2sZwVs8Io1THKkt
yloAeH9iCe+ZgK5NCi68Tx/TSqm6i9JA7NZFjxJ0V3ECy617n1KQ7XYOUPI60Rjv
Wt4mcsRQkJEYiW84XdXxPwrIL+awVkeD5ChOicEvAVh4msG39Q/qztD/tSPAgjQ6
dbv9C1B5VdueP2zw9ZWum+4mqhfEshuFon+vybklFNccKrfbamw8n8b23rwGihsZ
9/opDopJVTGebH6UlDENXLTZdycXUbXntg7Zl6o/RCef0cARW5I1ACdKGaNAn+Su
eLjRF2u95LIV2wQW3L0Off0s2IXPsQRMjVEO40LMiMVk1bNzaChsMS62hDojzpUg
2Kc7ooVH+PmG5cNQNcTcr/EDsy++kWiJU9ia0TLymbVclqG/HHKakphcR4I60sPr
5Jr0iL6Equ4GIHfbzW5DqmuA+sXABqo1LakZjnFzoVwewDvG3KacHl8LZwrHw2tN
9vSfOj2b7bZqNSMQZNyq6T2PHlIhBSr+lSXG0Dkw+78ixX9u0XLHiPLWJv76h4bp
JrI8sypgPuiss3AuzRGiuADSNT/oCij3d+MqY+tGHd6ITesYr/saZJS+hMmm5293
oPutgMd8wcJXhkKrHU00sMQXycMi6YVaG0Oxr8IJi3/sh0NqRt7c8eWzXDZA9NBv
W7pXtP3ZxcsYwOc2ECcwPOLjy52Bb2vbNSQVEFg3Tf2VdAUN2a+/UPhdTwniO8oF
6qWi8n31rrbhnPFid+PXChPtJPmR2HDwKIoFUZ/t2gSFtFLT+VmKTXGi1wEjF158
x/CjWk5/m1Q0pAjH9zkFldqm0OtRtDKmyt1zVFQqExAxvka9VZ17U603Eh9UVSuA
f2jC2D+s/lCsddUptv3drFxG+uEyyNN09q+BYYggfgpgTthUCr9OQgujbDYlfnvT
e3WetV37lYfMczXnS+t6SQcIO7+UHbg3oJp3tX5osibYGTN7U8rIxv8cYmpkWzGS
Egjte8ru1x/nDbiFq90R21TSHY5zhRmK8z78/Nx2O2jKp/tmDrqMrUbAEbymUDIC
FexSIKBi8aSkOz3VNhCmaGlkYWZwQppAGDE9oLjyu3JGPHmyp5bDoMrHHKk03qlE
DrFBiGfYyjedjXi0Dg2k+FhF1aTXLe3U+7DfrhVNCH7BGO9GBcgi/gtObpRXbelw
J2326uFw8Cgt9oD7zhNWkAyH1nTtAIkqUrb4KManZNZ/1fncrYtTjDo27ARVMeKP
smG37gKzSI4RwmQ+OnXxnedvvTVmhRAyj9Et2eAavIxTDWmdBh32Jl1Mit631UGM
If9cF8ze6SiPOLf9muaExIlVcVlmwDLblKHj+aP6e0I4MC825IFm6uUUS942gDYu
kCBw/xZsUu9dKNZWPvGnOxj1F9Opz14EahYvmACGLBF+BJq7SLRVffznJ+Fn8MmS
2pjkA7K6gUgRwaeCXgEkQQq5SWYYxGGAtsE0XxLvCstoqEhx362p4Qfdtqw9zj7K
3cZA10tL7zNV15Uvms086/ifmxUVodlLkofnCSPYmiXFF4ar9Aex6PGXu9vd4zMH
lqw55IZMKxgXev9nc1QTZBc0mmUMHdQTzx5yeGA2zzDFkWAP645JflMWi0Pfimkx
7dK0pJVHw83weKQsOQT0vbyNj0gjeGlHn5SBmRLFguyzRKmJ3w43jQcB/PMdV5kF
8pm3CAQQDNPMv6Ua85yP/KpTD6ks8us03mdwjI8rPQqNjd5oQ6Pn+1k21CIxeL5v
agaX+SAsJbPjyM6Vu04nOm4PIf3iIpzwKVMcJ7mXB8kH6HB3lPzSC7P2gR2W8vyE
0RqjmtVtJIKkoD1+s8wfqRsPV22JQUU6o7gAHf43CBczRA3sphMdVYPGIWCWPpjV
XkG1rV0i03EMQ6mTSdF+3gcrJoM31HanHYPXPF224y+Da8dhkTbq7BNCw1n36Khf
GdagKzr0ySAgBQ9b2KHbMKIgLAMNPmo5OUkJA0ydeECj9jS6RUzljHmZtRcV8VNQ
tOFUpA6vAUL6q8ZN1h4ZXiLRFF9lKKvTHrb5bEFFoR3my9egea6xaMNNzsdaJuvJ
0neyppuN4+ucWcODGI9hV356pf6YRBSjpBila+uprHuPax5yeJUJYhz8F3vdKWOo
pduISpqubU5He0s4WyFA1ZgXJqCEn/BpyxlIt5/XCTLWFgLYPav7cwwtsN07xFci
Hi4ZPAlELqTT/i4b8B+OKAsCpPLhpMBFnn6s6JwMU6BCEqtP6qJdPj5ZB9ZNFvkt
YNSBZjzkmu+hcECJGHbpMkEBahV3LJrH4y9wc8z5A8OI87x+QI5N1TgeO1E7Wt0U
d5GgnPiw83YIW2pamM+c174YlxmVascQi5lTk2ACjGPAMhEH8BLCG3nJOV877Mig
yksouKzmr9hqxUiEyRKaZeZ+SvuZm376+JfaNl4L+/8anhuBnU45FVbpPu+V1St9
zHApC5ZW4UV0TDdfAnwJxlRrK7EEr+zmz6jRhn47ptmGFk/51Pe/ocEsD3eJnOwB
esoK2xV2xinvDSHyb3+MO4LlLYiAkvLZ+T1mK6JHKlJFUt0rG0JZMtkApBZzmEQ+
oUMT45nET/hNSHGyc4p3CHJBUE0G6lr4gU6KicLxiCGjoEUfrvi8REXJMugD+5k6
vRumYXZZmvZY4rDrGXpMZFPnYLJCgUPpTM/mVP2YCBjeGukaqOKnwIoO+ICTMMst
ivZapqGpVo/h0vH+Xt+Rf7VtnealcI4TQ4u1ez5Uguqibvph9iCyHhWWbxG0BITX
Ccfi/FAiYUZWGX4GMk+e1ZuHLYuCOI8/FrubiEexXGL3oVVMilKDdsb/TWbqFNF4
teMzdBS1j3++CyptOStAWV1u2GBQTkho/Kp08QNF8a1hKRfNxkTVvhA9pMp0mlJ7
oqSMoOWCokoKVYjtqKt8jb98/mrVPPUQpKQPIueVP7BD7NQavmNqFxCToULu5CNA
NFnApcnK8azeAZKwUbcPVmNonmRiOrpschHR3P9qOwR2UAZsAnxP3jnblvb9MW2e
SKwvI9CY7K7oTUVQ+bborD+lZHRLuUpDH3NZ+OU9iwNBhOD4dutvXrXw5xwlJySs
Re2/dyEtwZyT83wTKQ+/0gK31hoLbvAUChNY9333PNhnD4yNxwLAW63F39NN5CHS
MoZV3kmf6W0NjAIh/F7ajCNxzMvIeYILNLqR/+myFs6WBLh5Z8gPd5yrf15sp7jv
nzkyZIFtFykyFVd835aDyh1UfIAu9YcwyeTsnrEMlLXA0P/WGRIdlJtLeOOXqWBu
1p16zvPmSESybFZe8KrUP68qNVdi+UoAK9WY3AtvgAZkmrhMoSoqXWUNn8GJXBPw
viUXSDtGNV2YyIEQd6cHgbJpjz1R7YZzc7NyXkK0Ls6g1f0iGcFYNP3truVXzuN1
4P9qqnTEXtYtuVUV20u6uXeVTIRSbkDrAqfHSInRvTwVbvYDkhmM8ZC9Sedbl2yW
JuPdOGFB0iggPTu7T0XaBPQJzEK4WdaImsgI2Tc/RgqcDFjE7ymlsb7bH0uAIZGe
3xoe7NqbbZGpsvgmGro78kUfr9b/dNvWCSW6I/JTtUiYhnwVRMSHboqTUyCUZf7V
1EvlZHilkOdjeEnCe/m1/Odtb2JJdlAMdTz2yBgVhk4WC/Q2sJTW0+x0XrNGz6mE
Yqow7WckDj4hIm+nFpPhXLcPphbjtK8VpzKx/Qf+EHMncPd8OzbZP33g5UHAlVy6
gObznskvRyg3BdkxLOCbLwUwmLqvE+V2/9SryupxHI+AZTBaTYfKlL6ON5D53Gpp
6ty6HjIPchrRZ9+skznDtgmHxhKYINW7C2m4Qkwy673goFYy8E2P0oftf0Bz/ybU
qrbQ3rh0TE4/YgWUeyOXgvF60PzK2sL3m4cCqju2SVLdGFaeSelvyX5QrFd8//rj
tSFJvMvjcZLFIqEQqEUa1rBSVxwYwVP7W5t9dUJoNPOVQDztGgHr6gva6qU0Uyzv
A6dWC7LusaVKzBVW8zWquHhorV91ExUH9YA8DdXrSkFDf73CpiTuNHgr+ryW46aq
i13cnp/5K7FIng6GtMhqMoMqLiu3l3w7QzrWlYw094xHQ+/2uAmU3B1aT2pTwoat
l8whOAQEiuhLUTKm1yz5JCrWqqRH9xlY2pNZJ1VKhsJxUO4w2Hno6AHraPUdgpw0
f4FrfrGvAg8qoWRhB/yXov3E77SGhqhc6VudvDohMgYvfxegVfzwbvV30t51MHOi
tqYc0hSj9YIGDpSEmQbye00z4YerwGymPkk12bntJw1M6RZv5fzEWPWgpV3oXgpK
Yx/6pjOi9fFi0suXHueFbpLxAiINo0hBDGcK+fkxQfzBdzQkL6ONzHDaId/IsJrs
XinLpxrKl6La9nl94UfuTcGqah2iv9CGv5GEunqkapHL+eu9yC2DFLAyo9vXKCaS
iW/1HR8bNZvYrfShiUX90cz49LnsswAzFoWl9WEN7uYXzjHpn74HHq+n3V9dE19B
+cCs8EYRVfXtrovtF+Yui85shBfXNZEiBfacLRUv+Lg/EkznoucRxo9TO5N1WveV
FWHz+FxgIktqDJ77c8MeeYLsDh43tCSCl8WQ5wiCptetxn+CSgy0u3V1kBOynY88
wWW0RZA3+0L3LHpG4xXLLCl7/uw1abwfdmyqew7tqmRlkbGtrnNM+aGay1/AOFmT
XzSm2Z1kFlv3o/TEruGgxTzwLzmgrs/ckzTt11wfcnwkkWVMYjVQMgThXIiJFoK0
fsgukeg5Dt8rbg0fGHF/7ebr5ATviVkPrWYYQO3/oLkqWR+ItNXhpUu6k6cDxN79
zN6K9uV58nXhmCqUKIVUdvVFOMpSmGu1CgoXHz8a5UklhdOa88rHrM8iom0vq8Wo
IpBbTK+RSUKQF8Tl1d3I1g24X3Df6RWrK7AVy1SyECf+BTCTZ9tBzoZfxJr2fZtx
+tT0xTovxxuJNLvXkgl/JHPv+S2qQ3h5eFR8MY2kEpMyAYFGAqmM7V8EhjPKWKWh
+M3bzaGAtz0oK9PSdSTMRMnvl6ccsfjaDK97lQ/hiQWBDNoS4tqZZBMe/yj9A2DG
61lW8/UsmuDZoNdP97pUW9dlih7ZncVxkCaAgGNr8InhA0qRVd0HAmKxlFVSoWHa
wqVBGKSOyQZe4rkRBHQveUv0HYjgelt6AiVtNewAo4IsZzIhf0sHsabm0BhO0JoQ
XC6tM0VpilYf6YP7ioxhYhh2TVSptomG+Ou+qF86hTqhrRLcXHyruHWOE4X4ToTB
EEEu9wLUSE+jb7u9+7LzMrMv89xaqgcJqxZAdca04t027TtQC7KG6UhshcPxjnIo
0SZFv6iCtusqOP6R/oJazgCg+Z/dF9ohbz8mH3wRYdTSlOn2F0rq6LRjY2T8/aBV
T43cVf62HpAkDo8S6f2wEOp+dAgZiTj4L9PU7CZkrEAYEYk1dSm6b0q82zpenVhD
lE75ZKA0OaqQhuGcBPfujWYySrFft6WvZGvYHTCTYoyOuVM5B2IsO2WRR7RwbHB+
C2A6gczv/FhSuV5vrD2OG+7GZogmQOi1+b5lnIzOl0YQkKuACyQy9ksA4uynrTEm
J0nrQN8FlpW//Gcghb3HE3QT+Ni+AlHvlWfIue7xulgia5osSC6V06fUu2Cgeuci
OeBjTqBjdMykg8B80eURig5wCdIQRatrTkcQhMVhwtuzPAHXCFkaDTNB2JBbUoDe
qq57Ww/aR0V2V/3RkhlQzEL6ENrBcOBFOx3ZbGPui8i6LsiWD1nEkGkHcHQEqcwx
3kP+L4MtBfboq+uMZMm8CYU6BquNFkWsTm9ZJdQ1lJVg8eIhyugy6O9QJ5+TdUxd
8QK7wwWaZ61vhBJjbJ2Rp003+m2ORr4aPJnMM/E7sipKu2J9qosNoqpgf6jxVnzc
5xy6yac1HT5I9loI3NygA33nsNAejU68P0CPC2vOAYfST8Gkf7en13kCqIQ8MACm
ueJheF47Aq5zT4ULngrrEHB39rDYPRktZTLAAQxzxJFjV7KrY2/K2CivHCquu29g
rQG6Q0fR8sTZkuFklM2T8O+gjQRH1YR1fs3E9rp2OKGTUr/hn9IuoO/1hE4tKTFd
japdyZ1eVGYEYDILFdyHvZFChObTcWFTnAfm/3naM4VmUTR1ZYERl7od/UgAA8AX
pe9FBsHrKHefCH/8l16nLuVqaLURosTW2uey7m9L2FqWDVnjN3Xj0MVZ4OFdEfP8
5Kf9T+te3HBti243aftaa+gPPJOtDnQDdpV5D457snk6cztE5Uv7KiY9/cNmczpJ
vbgxoffa46Ifbcc9talNV2FPxWOKODe6gQMjqc089s2Z+lbFWDQMoxKQUF9aBzHE
FnKeVHbicwGaqAIUy8A2aUSglOSAukdpDNSsdohd5VoY24EczC+WZxpyb0E5cYpp
H6pYPByRiP8IPceDzh2LFpSPiN5ih14v3bJb8dAxOPvv2YH6ephE32iy3mnQ4ItK
5KkUsshhkPNl+wcDMyZfpee9JEwmYPUQW2RKKKw7V9jDotGeHMV00NnfLLGdKlyi
3QjYFC2sBrr/VVC5pL+cJbt3d5U7BL9JYfrN/TpleawogI39TUoyzIrmf4hBcwOS
ipPH8uAymGiHRdpmILqnLEXrFwjsxlRwMomLIa7U6FPNFxCDBTx5IFyrSqVO2XTx
aH2jR2J5cNlyk6Sec6WsKZ+HisY/Hu29cbIrpyimCRBOqL0fxMRvhC9YkOMEqwXO
+fHccm64VE2iyJU2EVVUxKea2FAY0OeLduG4wz3dMeVGVUfmma2JSxBkj7o2Pz3O
cXcVYCb+pjTLcKvDRCftZE5st6dPuWEykgxfPwyHAce56oNWZgOXwhF3Ujbl+AAP
2mHZcGRlMvNnxxqvHVu4UA1u5df01+w1dPsM83cD7JtZIZP02G6GurH+ER87/KNb
6b5ioZOnxKlrx1aNBfmQ8BadRE5GQKaTmFrPKFA37c/VJOLjETrjbUEmqkTo5jX5
S6miwYRdGBz7a0RP3lFK0o7idvgpl5D+vuhEr2dKefwcStPvWWsVcUmnECtxcAf3
ZuAKDG48Gv+m4d8psd43Ls5AkTHH0RwQyBmoWQSqra9BckmfiXm4WLZj4aoTtlgk
nwFoBk6PtEFyId88CmoR5p3xNKbEphDyZmF/RBXdAMjj8ceASLGAPAlIbXX7GlNs
PJZ+T3e5eTsMuGnmJRKgi1/d1eLc9w60q0LA3uJOzILGqE+/rU7ylRwA+44K/5ac
axFPwF+bq4UWsTJ8urMgTWcddv0rgaOTiGEA65Mf6e3m5+8VVoMtmup6WUA0EogR
5i11y39TL3e5T/WQytudX0dvrZMU1hOfpoTyXrhz9V77kfRO46oD3mmsie0W3w9G
/PrKVtj7iSaG2sekMrurTTW70O4X10s/Sv+mBLGPnI2Th1juHDewhB6qI/DtUEaa
vy8nt2SvgJmEOgORMn0hoqe9NyBy9jbcJdryhSSwEIJsZ/1l3KbrUMNCnRC5SDyX
LKVarvCD4By/e/WUdjmEFZrMUFVVmE/ejaTHpoKxDipBwH2xMXirnpBNsMe4DbX6
2C+qBFWjb86EcUIkMqB1QayRS32uz2UwJ62HRXpnogCmGdq9MFldTrdTeehvBKvG
juBc+rQ/EezoVeVgrqZ0pa7MAbsKCRS01aYa7TBbuhtlUFJXe06WqN7iIRVdgHBW
6diuIM+9v4b15zyNoaJV9EDJRKsZqOVH+XG9QPejL9IsqQyUkmNJuL5ebaKJ1Xqg
EeC+4Q4ielEFgKwUqLRRuhK+eHEYISB6qvxdMNHxX6/HW52M4dPFanlHFQ9C7fog
aGf6EBX2FIzatASxZv+664ySaRExsulH75Qa9rxx/elO1FSZrK4tOHZEMwkplPgw
YKoLHKJ9L3ssDhDKVcI1u9CurWDXTU/DoEnT2CTSTMULbcpPcbFbvF+b/XFastt4
726Mkg+GdruDgBJQ2Hmf+T/o16Qs6i3QEv74Uk0dPrhGWY4tDV4g6628yz8eIVf4
0wGokQNBlXZDFkVuPrcdEejZhPe0+TQ2NugaPNxlgfATN9ABtv8j51g6cRs6ME1n
Pi6unLymlZ+pA1YwnP8C3VygwYhbnjq0irI9qkwOhq7GqdiOFa9dx3OBSAzZFCmo
KzoHKQIREcxK9OnRSpypUKK9CcLd7GVRmAwxQtwzMijk8lXK2nKJGSyjd+sZ37oI
+XDgbzkaKbTHc1UVXYIFEbs+H/gik42FtggcAsaiTnSZ+M/HHZvjBVBnEsry07l6
zvR6L4wXRcGusmlPZ2Mf25NDBc7YAVKhdCXSpjQUCVLGA4Iw55kNzeagISAs5mno
ZL86kVAQqeP+9NiLf65AxCuqfKtxOtBOeqJc0VeiPUF6xsKLkLcACSfTn4oGiXnh
Bun21uf9/EX+blzcz2d3NcYnONp9dcSiVu6sOQUqZk1wsJE7rSNNrwhFL503AKUg
OgQEoEwRvVFdYk954NB5N8dqWKsPlZekg3DDLdLORxRzkSHo33kFR+yWwe5JWOY0
cdDCOF2NJ1A951gSgOyJSI41nBlhNO9cxNr9eeOqgk4fWoql3CXhb5sh5ETyI6/4
ssMf8OnW7d7oCz3vPtJriyUM23pj11oA1lvk0vY7e3GjEaQxdYDsBpYWL7gHazkX
211JEzjhWWdHIpts4aTv54X7CaA1UPOhGPKu0IsLjGu8M4GoeJIoHR5nYvlk2yKt
Ao+z3fTqymM3Ko1XpTpUEzPgPDOC5PB22WHxNctBZaCDQk9GcEUly7jfn7pYEdMN
/fRye8kAYxYcNtkMoYQJvCQvyHj4lh+UeHAHGJk5ej3bs8gEr29KoiZ2v3rcpLZ0
1vYtDVlmj6LiFX8//nk3cPaMD4wzwuVHYmIMYrKY2N5S9mLxOG24xefahokx2n/0
ico0N/C1ip61Z0snX6P01I5O1VGISdqBpmS+ZCwTtUF5fLmdQgaPTGeVPNxJQ36N
nDbutmN1udav3/DkJ4uLS7ZnuQRRd7H+PDhAWN3E9TAC91A600DN7KVAJ0Cocwib
XqxADQQ5qL8rErejSLmoYXGiQY7QhiDgjQT413al2MMhGjaxxg8Ms8xuFnY7z6m9
`protect end_protected
