`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
rsiD6tALCqmGpggWuk0CLtKfbLEkgRopDqgJgqhLJGbs4p7Xl0ET16fjtkfkcLPo
E800aCMYKmZ3keyzq91DESXNe1Kewr1Pdk6Y7Xn71uKbTyySKu4U3rYdF4yvsFR6
o9ZAc6EszxjlE4z5JV6dVoY4kg8aUaBTQaZNaRRWeaQAK5m/BVH0L5jnlaD6Tf6H
A70TIgnU8eBewYWScW0a2dXEHS0QWu8PsKX+gCxdtAXwp5xPYxAzSr2RyXT0tWc5
tkolsJMhLVw5QOCetaCj0eDvlOGMfa5tJ5Z0/Kdbx0dMy/jcUCoca+JoknO6CvVc
hjQqHL/W6CMZkJMnUNBmVw==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I45kUa06z2aq1mAyrit+/H8gjbsuzz8hOJRN5cha+WW8m/sjeOeYB1qnCwqbZfda
iCMBMJoQ9o/r3J7KlkRQh/z3kjS8hDeMDErcya//raWlQ1d7L0BchZHoITfFAwXg
RMyPnfS+vfMnagTVTbADI448VnMKKL0dBH38DSfiTQA=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10128 )
`protect data_block
xa7J+Gd2SQv+hhDB9azZULJwWwddnk2hfvpEem1nhd5eplagCqGB844F9sUkyDWi
4u18LiR5yPjrqzyY7YtGByWneacki0Pic11bXLll6goCONlBR0yA/ve8RDFZ6BiP
0lBpGYOP3r94ATej48EoJ8XVAkqicHozpM8BdCuSVHBB/nJfl4DXlDRey7IdIWQr
2kNiBV0BYaHqzpTGwslGak6KIxcE2fKesX0WcMa6WGq2Qjl9uREEzTFJUPd9+JUc
WAGiQDWUKs7mjLrnt/jqDRoCu2amJQt5kmCnXei7gA4BBDp1ArMBMwlAoayIn6UD
4Q+Z4DQ0x/aY0uB+dD7YobJS4gX0M/tgkc9DutKSAu0OMfOwUXXgBiRLtznVkZHA
OsJwG8OaiVln5maeq9T2YVXlxh4SuCcpf3yIoucdqb0zh69d5H9N+uSm9gn5yTRq
3dIk2Ew5vU4oIJsdSaZkVOdJiljKUqNTgeO9NtAmZdeOufJguqpQ4PdadZF/y/qn
PH9qerVmOOMtE8QpKtWbdc8eWQlsemXErLDq7CHuVJlx8hg/ScNNN4kCO1c/JwxJ
x8PIh4RZTtdb3m2LLgWJRb56PZOHM5xzXCk1rWVk2bFNVQ4wqM2VN00NTxYsmurs
kc3fG9oMFdjDvXBigi6f/IONbEhAF4aNndmVEThWnKE5X4jg4eNXOz6a63XScfH0
kbgJ76ILLfgnBPYXmg33cLDuEG5kzTusfwf3o/vwKhltF/+/qeNrO3eMzakjHVnH
1fmy29K0NgZW29v2dazhinIyoKoPHlGjoJLPnwsjF5AAVYvBOmfMgZRO7BVpwZca
ZSz8pAMiPGuWqm7tTUSt39IdJL2xebht/LoYA3iE+/U4NC80rQLWYlp8i1Fl9WnL
LxqgalYyLUjnNgp0/y/E5Wjd+RrJRdnK3/M2TYr3R9UAd9AZMcltrO/EKfImMgHr
8wMpj8Ga2Aa2GcnNnA/4TbQSYQz08a80mddjySfcpyEO7LAnRrT6oWvuICy1s8hZ
cuuG417ZJ4G7L+eQsVffW/xbCwF6DSn/lOVZ9GUGVWeCvuQvhKzq70vCez+XsCNm
LuN0GxG0Q0FoklCbvv3MCdMQBna/U1aczKBlS/isshSLqCbeXZJ5A7BwqAFmtSlL
y3QuEpXrXDI+NgYXlops80+5/MbZNAAoy0pjJVl4sFRr7wT5j6e80W53IlMjvimO
AIAS+Bcc+ypEz5uprr/pt4jJQeeE4Fgugry+lIxGw6RUh15O3rSdzOIq6OCXh0gX
Y9Ss45hhWopUVj3lYD/BeChJpmg8AQAWQV+ojrgo2YPG7Y5jxviurP40s5Ak2MCX
4oOZlUFsRsaeb5z1u3I030sMKXZcx6n5h0vShQWcYc6cfWkXX/zyjbo/8WpWk/YC
aXNGHoM7U9va5J7TWjJVqr/HkiVacdVZMiRxs0E+fJx6kxkUVaok9IkLq/tnb/mQ
wAeiqeXasJlAKSd0jGq22XGTfI26wh3DBtr9I/K5vG5Y0uHD66uxpHDURPeJn6im
rqribP4O1ogwZoIvvO/iJ4EvK+Ieyenu6VC8a2fBrq7rdANsqU3Z9YNKzvaXc0wZ
AhjBPmuelR9EX+RDCXtLLTZtih78WARLQPrGzUYX5OgLj3EjZW3SP8plSckt67Uc
EMrrcichyU/CG/+kx6dwKG3jEZWBh54bkYYYqRVeyub+EK4cWbc4v9ugBCQCqg18
Mgk3bI47lCTgTB01yVlHjMLGOT1PUz5dopKTwBTwJ2DGcPMuizibAiV7hOYgvIND
jap+TEBeyE34bpUN1jWGambawDSYRw+106tCNYAkUHGMldsn1rHitr0KaO6WBybC
USjjReXFT+6CrDAZIrQYY5QQMikS4CBI1/ksg2ayuS+kGlMYDS6LR2NVXlBQZ/PN
2tkr/rjdG3WnflrZ7Umy2qR+a6wObWPFOBPrSxNRJDyQwzpBthd6xf8XTPrGbBoC
HlAsTzq9TiE8x8xBR5F6Rbcuf+VsXtcg0+KOWCTJrKNYDv5l/sLQEQbcsEu+CzGL
mw4bHc4omGe7wj2/ealuqsdj5VpcEMrPvFP1XNRfD2lUHHO8BanglnLyOmGfqr4b
MdhPaP7oN3ILeX+nl7hBzamoFy26NfqyClSoxUuGNZfT0VEHSr48IFznH/cy4Uae
61+1daVTjktY6oM7Kxm2J/qX3cmjX1h+lLOC++GwsdbRXg5/Ek5y6/081RzhA3c9
NznQ4UbqcZi0zbqgrIlwaYP2LN0LvJVfkS695pqSEgrkv2aMJJc3N9GGdTrFe715
H9y1c3Lgeb+GCz0l8ZO50jNx3YttXiqLCgya+ZHYCJZphR2+5zIIWTz00VqzmHjo
zQXiNWL4oUChzttb5xZdj9odf6H2CH+bninyRAD3zD1c7uYxeDZF9Dwf0a3p48+r
SkT22n36EjDOzpa0Md2EHTfeqf1fOQuKdSDVR8uDxkyEeoWwSnQkSvxGZoFBahbp
V5XsMft912lCqKXKvNM8tmuGchEepisC2f1vxecQyaffogZsHd/VJ5n7rdXKOmvM
ouAGILpxnjGSUiwow5HB8oSIVGaqcH4bjALJfume8DYOenY+tDGuzd4eososIFUu
B8AMhNlu0yQCemh6Tho6TCM3QwGkVxszAolKf03FlxaAZnfBy17K7hO8hBTX7g9w
LDox7m+l8VOfbBatWoxhMxQRSK2QuHNeSzGJywAJYJfhuP02ZFM6eHanRiphtLHs
zAUSi/kmTsRGNbYZipm502Vo5MzNdC9mCoGQDo+a+iCUyMWYENdFNoANgcm8KflI
sO7PNvPVn5QAHeQiqZOMfB57AlDkw/PjPHyOy4TNuIy/IXwd2l6ngtsIjME/Qqu1
ZX17IeqwZhtXsclimgDxHGlnTVL4+Arczpod2BHa0cL6TCCaKyhw7hJk07EgLer6
RFKKMlufqo7YSxE08Kb5llw5YDN0J9cnulImih4XvV8dMsDHAfRWFn3t5i2qk/6u
dhm3BynEsnFlVlFPeQbwLvgJU0MgwFM+WWSCjhC1EoVQQhXWJcuKxg7rY/oBYQvj
8xIs+TNNGZUySQYSbzK+Dk/ZADfcfon8YXFJF6QVtZJecagQqCqxiA79QQheH8Ql
abWbYGndMDpjE1T3sInCSP4zE87nxdbIY+qgNgUeP2DxRMMJbzOciZboQZh+aqiS
/nZMwiUCeFtM73qVk0IG47XLz+0dCpcNJfFtCOVO/1SKiwWhIvH7UtfxDq6L9gZN
3e9DA2GApX0VwfwCfGWZDwLc173sglBbD12n3ea7GuJInRWLE4poo7kh7fR3767P
3UYZ8rAgD+wOdfzCpQkhyZORgK+nZiVksSo829HW+EjuxYjoX1CyZL2URpVbxX3r
1bffFty/GpGR5/JR6h0xq9Tw93NMV8GRavrrvV/fSVntYUXJtC4NEArog6Tb9Kqa
Rf8UOh9Qq5kfXc4WazfeNtsYVGWxnftxYj6FzNXuH0FB4gWIEXijjq1sdnzwvP5a
P5459w41VH5t3TNLooVGzj0qRsAgar3GrlX8iIOSIngJCeHqrwdJQN0G71darFtm
loI4NF7MCEq6qMLPPfPfuRHXpu0PwlB2fVTT1vwihxaunwLl47dwz2h5jYvGDwSG
rW2LPW9u0gu/UqZCPW+ZeRA+Mzotax2wL1bWKA0nEgAzFtlRfI0P9uHT3rTEzU9h
h1V3vM5jM96MHj8ulcXxxsiaHwhaT6O+xKyXhVv/vcVVeURrVfx+JFqk254leelL
l6kKdZLYMZZo69JBYua6Fzb5cph8Ey/OAEa/8A8sBtAr6xJylzcr8QxfepJSZ/e3
rcCnr0PFE3gem2i597d6vBklcewHSPjpkQbCtoGjI0+R8M5A7XEa9KI12fqe97J9
omVYwgV7pp2V0ypKp1Mt1QTq+IF1crkTx+cwb+12biRAnmyBOnX7jWoeu+oi/8eh
89FS+fyAibEUKWRV6YcCESQa1oOpEDu0V4Olz81QB4kWy/+qnzykYT5WaAEOy4WU
3TkOwrHofaWEj1Lv+m816ilGSENtSL+JMvz+Rc1JQBCr+/QmsSydsNOC2GoQ727T
5MjzqHPRdmBLJJ7Offe3za7TO7SIJhpJkpeZyUWeuIrGsaHjdlmhbWsHEsG3gtde
0ULonVxFx16JCSl38VBQ4nBzoeN0InvyPevQUm6lCYdwEadWWj+txcwsWu1zIGp5
Od1sto/hzFrS9fWyduZLBWDcc1fK5IcQoE2MF60CGTMHb7YDikwxbwxz17/cgxXD
xj6SMiMQXe0anSU/wJddquC1XReLGju+aAESJYHHgmCTta6FEc2TZ04KUDRNt6w1
UzDHC/LsakhRGwW4LZ6XoVtwaQuU+JAJjnNZ40oGnm9HN/ymMBgwJirkbt/zhDtt
xrWY6tkOs3W5ncBXO+CD5I9pKyrLzkN94Yw9vRmUbeoBI7agyNevTTUgvIkmLQCu
6+tmgi4mSCJFLbPO4C5sqYd14N9/MMyCmkiy1BTSjeGPirTiV1VCpNBnwI2bDbY4
vK03/HZJFYxsSk75U9lKBqW0lIbQbhjsFRFXgo+PQOkVsXrBXW+NFPV+5ZeSVoPD
kIqrCnaJpiPLrUqhLZcdW8DgutWnGX4vsOh9qG/kKW4Wq7f9a+dynqu6DO6uhAQi
77aqtl2pIbxwft4NPDR45hTgBCgQZTAXZkWBR5iXlW2S5mME+jtMuqyt66MzrolG
KZwoghwyzasaPOIw3wqcotsMYlcnXNOpcbYeaqha8j/aSblQuYGWcndOvhngQsfR
+LQy7ivnavVmlWel3utV1bpFFNo/swwaIpINPonHQFmY2csthdH/9Crdq9xy7ulg
2uLOmlD+tK3zoBIoiJ6X6+abCvyFNnz1BCFSGSxFj5y+sHmoyQds5zQ5z5Kz+myq
xRssbV8SSnawBgG8FXX3CixOLxwzDrrxHINglcMo0/b+pwP4tMJS3J2Sftf0PQRH
trOtCgJO2eVtRoVZ6N9Fx9gbW2IovXDfq7B+KpMnOAWyyMXL+yW35vZhO3zcCziZ
D9zNaFHCqpn+iT5kVUwZ6oP7wIbVtkrffBas5ac9lvXvH2ObZzaXgnQQfZGyuwrO
QTm1asXkSFoMjXEp/SdGyr3rGwKa7zEqtxv1ZpJ/cKwOJ/+q9TAG4fO0dBdZSkp9
WJ4SvlyMLtRhlzdAq6RTVPcMOvD0o6oSB31wLdJoINr6xIYrzkWw0xjubsf4A9J+
szquAgk1rd0r5Ya5uTg2TZUHVer37ecx9wQa0TpTBKv4wO5NrHln7bn29GaJNrjJ
SWsXo7iJx0/f98wwRJq28QCQJ6vPPJEquguDlpVagPxTHYkiUBOp2+Q19AuNegIt
wqQx0li0oQyqw4rmoOm7P6zeumaYW29yY+mpQsIplcBJoAj0bOiVVCotjkE4nbci
N8LrhQmgx5DoZNmdJYuwIuLrenoBlm1OSlUcX7UntiHlB2aJK6hyiAssppf3DTes
PjbrNZ1nYBSWfilYPd0qdKtUA0XFpG/ShM2PsdFhmYuwqqJrDF/xnnKmXz3v1Uxw
6kZGvfnFrXsuMiha9GNLSUufF7TkwKBriy0ugxvkvmh/4vU2vt3olS4uruaokKjd
61sClEY/s8il+oBKbzaDENuhXCjRH8Ld/Y7uIZ6lKWXXuhVZ4Z3j4jZ9Ma+0rQjG
W+w/o+hvOfqOyx9xgLJ3vFAIvSY7OymCjXpnjcJoZfQx+zzbRftKzWrQgQzbSZwc
Zn+YpJRITl36Qjsa1Us47SUt4u7FnpyPABvf2RhX2NbrVwsjgiGOG8qMuJnUmKTT
R69TuDq4k8yVGmMX6XaaKcqITeiQud2DZkrTVyR6SuMRKT0jL7G8AgjK7ekv3eTw
5Dvc5b2KXs5hBDvolxIf7BpqeqEjrcSWqFixKinERzFTN8PUcGIsMblmPHqQu+0D
3qWgSBxej6A8xxDVZKESHpVS1wnCx2LKBT6YKCbHj7m+J3zXaakUyvFZkS30g8b4
q3s3/wx3Sa79oM9D94xThNb5v2l7jNiopZ30HAjfDY2Q2MkcjFF7Y/HI068CKith
PzC/tpV7R3xKVM458IdrtVg0+8PGIcXJorUFlZKmhLrzUK2EKkLSoxlEfFcAN5mH
eZEcMvJbQUSfBjScP1IEXVEvebdz+AMstH1l/Ge1zpyCmGbEKwhrF917/xtgMqku
d31PAyGHrxeljYPBI4OZ8Devx5Scl/PCgvGUVvPCyQdpnZvLsn3Kwp6rFH8X8v1x
dJEvlFooB7Aroh4MF+vkOdEjWoEmCdZGAlOKnYkoSQ/2sLHdqIuaL/Fs36Nd7I40
x3TxztvuO4ERVa/+ckkw9AFPAWaBIQiRi9iOP9QgMBi/Q+uf+8Lc+UWxFSWsf7gz
wT1Wt8miRpxd8ZzLGPG1jfvxpSAlaxBtkvh4gFwWGI+Aeuuar/T97cvF5wCpIv0K
vJ0RLpUu7KokctxQLuC3tiV/n+iIHWZDB3fEvBIgoJaiVh8X6q91darritzdX7jJ
rflRi4LO6sHf5llFG7QsD9bkHg3q7gQZfQHKqkK3I6oSw1Zr7FTbXqiFat1TqQAO
G3kUN/OxrLffcq2rztFxjIHIhxTys/makg362T/bqCjHZGALZjMMofVWzFPHHVM+
CmVgAmkuPJd2bHhan9iIqFzgGvrBr2WiXAg9bgjX0aHdhFWvl28PMOJhkl9H6ftW
Z3POp/KR05iGPi4cBOhh8yf5aRA4K7p0+U+w5f1uwHxnnCAzUB329USkVlQC7YLr
pHQUYmYrEpumMzY27LsZHH3n/QWBgl8/2vdmFueXPleMXTkyEd7SXKpxFxwtta+l
wJs/dQzYqTF2q63sPk7OxqRady293nF5frpgRm3zJ/blRMV9uDsnqvmeCHjrQJne
KQbANtuI2fainzwyUA3hkIP1rnur3FctHTIUgGx+dLsEUGjTUxoem5+0FwCu8QcE
vzgUj7x9sGJk+B1OMkI/h2M+r5Qt4TJnAhnGhuTk+oV5i6rGl9Ro1lWiFRbS/leU
junVEQEAMGUvYKiAwAU7JGmLKAl/lTuwrSWB2Ol7mfLjMd9TP3JeGLIpLQCm/ga9
khbLi+WBwxCcXVwV3lP+h1TbYNslxHp/zQaf1nbPp5QRuvZzKfWEiWEJZpj9iRb2
dz0LVByUwjhcFixqJucIOpXMYlzA4aP3mdtcy7+rPeBm83eQlaGHoXP+a7kwYdGy
T+c040zZuZPk3aWEIldukniATsAK1/bEpy2KUG2E7k8RwHnNZcE6fB+yrubUsDM7
3YejSASITDGUQBjhgbi/yFXnWqnCXkOamR3QBo/AU6ZA/y/gDqMcoL66u1062HtW
E1QaIPeRsz8TEodxg3CQE/j2o5sBkAmHLCKyIS49MsSDCaHj13jcbDFofIi0P9Cn
hYYWxItr+1iVHJ5w/jXnEDHulp9CUZSck0vo2mRFgZ37B0J7/8Af6CNIJuyxKirD
1ywmbPjkLZWa/3hGOIa92Jy2VrG+MkZoeMOqDNwEUtL9/03cCGuxdqQU7QdpeBdG
83+4mDHQWK75N+Yz1/q5wZAbATlMKGl91NregFnJbwzQ/+fWrwPI7muIzqRoYqU1
5HsBEb+FzGWJ+0qBd+SAveCxeD1Od38nhUVVibfXzoJumBqOcK12B5RTXBNvonjw
d6MaTa0ZeqQ8UiCGdA1N9pZYYLKKlIXFOh+7TqUWoMx3i1pvtrk1rFCdwAP2MFAZ
ardpa7+rD6ya/aAstumfZ0Qe4rDrCHy51f4TU+pdx3brSAX0mM8M2cChVUnnHr2d
B5iyObU9inYUa3+aeCiQVsnJEX+XQ+Qt4uZtAfaKPdCWwSClaOaCj3AMKQeXVdmI
J2nwjaLn/voghMZUjcxJarIVPMvAheMBL6nMjYmN7rBe+IAFAawpQdGSfRtfC5o1
+2rhJfi7p7IiPKmoadvHak6FJo/RIRc/pVq9ODH3yMp8e3uOWLTEa+m6dIUqkKve
xQb13XKZvzkZAXn8KJ7yxhp52gm1nkqAKJ+IBkZ5mvhqVgVNzucYc+ym6e70DmQX
Y8BQlhrdZOJb+MVbZ2TMVyttPG7FRIDYKIQmA647BHVaFsDweOGpBRrISJRWFoFl
TkeVK69JEKeTU+gzmy0P55RDw+P2e8L4BwTbjzpCv+WrisUUuKc0zKOA8A+yJDNo
w5jRhjj3szIrNBfb8/uFbk/aM4wRIdPwBcuhPKT0amghqyYYfctiIAq6A++sUS0v
GEozvJzfNv5H9cSr/YZyiivrWcWbOrmhAMmZQlW3V1j3ksSN8rI7O31YetN4YSz/
TackM3BitMD0QS9f1aSbViNCHZKCwIs4ZsK0qek+e0Me4BZ4e7oy6Qs1wT6icq7w
QbsU1UkpWZ5DrVXD+aKVMYkSlB4G7KY7mwxOvcikz5PCcUOHuAYZxaEAFdPGMqGk
jTyxgAmFZ+yhjvwFbs0t92bV42dhN2SCzmHW1ma/eGSKmtvv4VYZUzNly959qcpK
3NDV79OX+PqSoV3aLnr+UB9j83nzphdjT0TeWD51ATYxWljEoaP6bgDgDN12Lu/v
KrSnRDPgwctvLmMYyuypUe532vuKAFbRDvZhaxSQc/aY+beZg8LyD+pYXDoDs7Tx
9CwbFbDkZhqItq2cYyuYRByZEiPYFHm3+daehfY+OENyL4mLcPB+ejf2+gJBFg0m
f/koi7ugJlKdowrVQKZQFY79JITJg6jj7u6kiynLqALacxgr+pN48zBkUXc6wV9R
A+3fcfwIo28h145oRrGy1Kduc06EGPkwnbF3AEHDaGpsFvaQuSTGfB3eyN5aiMu2
ujdoPpliB1C18Qaxn57+WTIldiY7rwOcDhcdz8w1l+zHiK8ryLV26jzMnjFfWATs
L884SZpgM04SwvoiUAFu1N3A0YQG91lZ08wExF2JmDamH4MK74TJASf9x3Ou3HNy
lDMevC3XCyL9yO10yBckr+frI/sj1rR3NUr+mQw+zRC9NRNMgYhbGnb3DOMQEEYA
vyJRPkDEXgCpsV4/1jEYlbMjEWPaSKf/DGZlRrzynaMiNkfAuOKiVHbhOZU6ZOvW
3Z7q1roPbMnGuxo23WHI76Ldv41G1Jc4XtwoDNQx8MnPXp6Ahzh4kM/bqKSEjTDI
AyQ2Y9IqaHNc6M4gKEeGW/01ff2wRWKQuCa41MSON+Nc4vC75UmmlzqhuUjUvw0j
0oGY0V7+BwQjFYDd0TTtHKZQ9CiA6wb7kEC6AQr6He/iKgB/YX6JBSNaMkzrvISs
jzCFC2BSliRT9ZQlJzt+J4w3Z0e17qk7upE8k3oE7kmoIBTtjENknzQLxcW1f9Rv
YT5MpV40j2102aqL6ETO13mUA/1L5h5lNreJbsKf/XzfRENC9m77DA3ejmEfcxCU
DBpO5cYbRk1zWzJRmR34Oo+YnhF+pHZUzHZw2rqruc6cAyuLerzQdSSiMXxp2LdU
LvgUNfKCH15X8FkDbln2j1N+taIs7SvkP+A3BKyHnKVZcGjkvWtlhPzt6sFFx9RT
tM8RnpbXsr0qR5rjrqp/LfI8bY+WLBxyF+viDF2KMJwwkCFOfzfGg7YKz4Evuigj
A4TE94FE1ER55/HXnVB+OIOvERZetmxjjyT7hFj2e2a1MJMdpIunQan3ZQofjQUN
Y9vMrAvZXxo/P1MWmhIWV4uiG88UQB8NpBYWEo9TK4iM41dNTnwEBEsgOj6KSdkw
pB72be3sb/hcEHEnRLt4uto5DRhkXTESfE4Lr5JSpOyKsoizAPMAOXCdvbgitSdD
bQJ3fVYJXQewk3gj/GjuWOZ2bFfqQvjk0aU48SJgsjhHA+eXF8WZyhQNCn0YOT6a
mHhrya03975VtvW31ONQor/uCvShSUfv/5eqH99SP7BHlIoeIKJ6XgWjjzRUf05a
N9zahvqehmoeykHphoGUiJ8XgR14ulMH3/1nWHX8auG0V1DszCJ9KJpHr9D4blXC
Rfw2Hu8RzOTC3U8OhR0e6tvL4oOnZzQVgn3L1Ew1aPXE8aCr4QxDyEN5SJ+CQXLa
hqlIDnWWjvy1R5IbjmyW7KFCJMkxanhM/Lxal8M66eZFlObiKNEyAimdiM2Pb4XC
PsBKfiLZdbfmEnCo/m+d2/9c3pO9Uo9dJkEE4E5rt3Yt+S3rUtxaTbNVhCTL8iHP
gWgY4h1/O7ZA3drpWXbsGeEt1/8tF7V2EI8ytcDFzV0iwTGNsFCWG0j3nt2g9LF8
jeH6LExSkcyaoWKMPz1M5iimn8GVS2xj0E3IYszeMtevCQABUN60eiS2SfUuTlps
To6QpIsDwFph7/Ic/YYsfCA/ftO34ApTNmwA6zDhSkvA+nDq6JJoBeI0Uij5keg8
NG7+d/oDsTsNL3LKnxmsprbcJ1zTjzm0vquSqQIwSV7wCPj3UZv+QVtMywqaEjAz
axCtJbItE0VS+MC3qVIydzzxuenRU7vnhSbY9/WU+Njk7VIIo1eLRU67Df9Bl7/F
KCyTn6V6GEhARkpGBWwMI1qGktr22/cn6KE9rt47ECXAXGkbkZgbEiroN+Qz2fpT
WOiO4Ll9keE1yVJbABHWpx5aOS8kFNzs5Z0UVQMaevN98peSk+rHZ/gtAlj4gUDp
NbonZgNNjbGD2j+7RYk+gRJfK2ZPC6mPrh3a6aXzkadw3xGqzHgqEHBrq7cXNP57
HfTgTtd+evG2NKMmsDPu7WBTOmLMckzwf81XlLTmdwP/AnHC/TjHAe6OX7YTOs0a
s6Rx/cvwSTzSibU4el4tp1ewNugsGJ+wfvgI1tv2KFR+Gy4L3I8VJZTdeH0o0mbj
1Gebb9xXTpXozB+WhWkkpA2NbQOjvNTOxaiUUSpepJvdKH97xwxCQ80l8Yxkkgbg
bRxafREGxZXaSOeuPBcTlBtR+6BpwC5sSKl4qGhjgtDpCi7YI0Pvusu4XeFBoNDH
TdLYH4gnsQFTSBfpHjPvobb3ji7vp5bXGv2UNQJgzWHtsJviV+iD1CTaLe6nwIXB
rs6aZ6Gd/hklj22iEziMfR5sBOFhdJKnOyB6zXQggH09ZZLMczjH55uC5ZUcbScO
0+mHtZowFWBn3fhbvKSaG60aHKc80709ZO7Km+pctI6bw4te+YYgCVI7KZ8tP2zY
x5JOmDXfUMghPeTbx6DYVpzdVfZ4svnyxWhtNa9H8P4ta7RhyN5pXgy/ynVj9fnZ
HL5zTL3KpS8yroaiz/VkAU2ugqdzv65cMDNRfuMitYnx/V67MF2QYfnOZntWYNWu
CMCmhAJ1Pac3WwmnFdop9s7OfEJbK+sS6iguSUzrAsY8+qpRn4hpZZJacoZK/5eD
yzrYXWGIirX/T1CgUyFrbKeh7AanGqXAM56vMlsFHjxtkqsbhmLngrzPHJ3NeJbo
Wkt1Lv3s+6JxW2zfRxdqFxZVx71RuotFNS/Vb+mvS1+X/LrWVofBZ1lgdpRTaSpf
Cq5NH8UCAYrXN+zbp3/NH7f4xKKl6Vq6Nhnilz5gg9P9MJNGT3TlSB//MGmIEWVe
6sAuQzyqVWawEjjgKi8ppgza1E6wMPGwnfVcoOMQK/hUCsSBsYv8dY+IuJ+8uoGi
rvBXC4VzS8Ig9NYlYaYY6ybPQDucR8axrKl7gROqaAHkAWXo6ZG0XSks98pzlf/O
onoy+4Mk8l45L2M+X8Ni5CaqJPNQKz3Eg/f6+qD+O1vG6hDN2g5u8lrJjGew28Gc
4OwLUvi8kQd1Tixm6NkILNEZZED3sXxIVDq00zKnduOJEiJ0qhHY/sfRnSKjrN3T
j4GGrW0vjVt4WFpeTvcgTTJ+zSl5Y3x0vwaosu3uFlywVtmPWbjVocd3YOARB3Bo
/Y0D4x5Y7NT/mhb9trAX1p3aHmided/CeEVEqIrGR8J+d1m7M6gHv3Y/OHEa8SDg
mdtMzEbhsvaH1E1COgEZ4kHoIiCtsQHemz25uIKU2+B8XLQ9QFW7fIp82kDEKwwh
3E35NILLkdpGq+238JlKYoO0SHBUFg5+h6h5kb4p6XU6fqi/xhF5OVSRaqZlcxA7
0aj+8PycnzbNvkcvmy44k0duivbTzySVvNTY4xxx8H7xPwQ9fvqRY3Bdhi1D8Z9Z
RUAAvdeXUYLd8cstbD96ZqSAX7ADriDJfKpPDkQGQRfskizpkzRYdTcEqbQU+o/v
HZ0GN+0ZgQ4GICxa5wwqHfgtyC1KvZzH9QhdNKpY1p52s2oJaG4kl9gcQFXNOyNb
aj2tfmGuatDvHohregNYhyLod+q7v/5XIuMNXfWeFqvHPGF7DnqBmwBIDvsLUvhL
X75RnUe8K6RPo1w03idmsfpYTEQCVJn8rGnwN2CMIXCiLvzEguqPGS4cqIVWpGEo
AKBkaIoj3HwxubgMBUfiSdyhdVZKe8/B0M+At/5V3jJIYOUBBqsQxmUeY5bGYcgI
JCVHTCmCWkcLS1qjfkvCbOEWxHj2Q9rXOiKCsci2NFljM6EYfYHQTVba2CMJLhuR
KOzbBN2KX6v4iGR+g0g8/WseK2bUAmcr2GiouE8Bb+299dvEW1s1y9YrSYgqYWmh
LCMJsNuRi1HB+MvADO1iJEZZ1DdqeT79KNr6FtTtApXZbKvqtzozTzgRctg0VhBk
QyHHe+wh5k8GkqsgEmnfSdesvJHgK924tgC+Jr0FtKvixV+eTxWEBbH3hZCrsg0p
oiM/eoAaX7+Qgz6ucMdhQLtJ56ullEoC3JUDfMMI4x/9Gy9h1tMVjSnf3S8t1OeS
FPs+Js4vgfer0FmALI0CIm69FaxWSTnlwAtfAX2wd2mVWfYaBT14o2BwBK9rPCWd
18I+H6KqTcoqH3pSEhZzEiK0qq4EoGnHVQaqy2MNLuk4KD5t7J/wkhVxdqMfGZ+8
YieoPd5DNX6ywtpQExmnULr81uE76H/ogRbVg+9dez+dJwd2T7/4W0v0SRC3qxvO
D9jAFfwbGMYqezfVHShXcW/Sf2EJBVPFAk4qAPsRM30YFpcKfdht2b+PYYnI1YJU
gIIdqlUK/MVwc+NznrFc4j6bARoyI+xukU7YeTAvxBi08oc0Y1JrcZpDROmzzYNf
FD8zOj0DHg8ulZ2wt6xJN0mASrNFWnRhf18+Lvv2qQm50WKHHN20ix7m9CrQvGtq
cOhr1G8G/UIgny4GOmtAp40kX4veaIxPY6FKJIp0S7ontSwU4uPPx35obBQ75Axz
FLSA04k7Ji6YHJ6JUB7XLuNn4DFE4gA1y+m3j03tTDRrk4c/q2l5q92lQSagrYmo
GvGMLMlz4Mm76BoWf8pg7OTkN2AysAZ8HX4WhTKwcz4QQJqq/k3nP1eCoa+j38AS
vZsfJ7BUydLkGjvbg28A0xTbr3eYQrAUGsDEcuWzlrYDnbMQwNR88yL22ncUofze
rn53t4Vru6rMvTQN2nTlgwsC9SwakmIqsksv2Aowo9YwFbdGGOkoITx2JTqsG5Y+
alSqY0MRpfyHAQWcPlKvBuC4oSBVALtGmSKXJr2btYiBOcoOlZHfLIRtIKSgl4mo
`protect end_protected
