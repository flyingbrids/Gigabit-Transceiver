`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
PfEDvyjgAKKbEdVhieyiuYzQ9l9WRQN5PoQ2tdkY3o8fAh2JsQW0xgsMdo2nWSk8
NmzQw8Bz2gWLCLKx3KUTAKxj8SnakS2IoqmthoiCHc1C83IlnAWl1s+zG5hpKsAf
rXIOMmlhUkQdS3MTeDcObyfTGbXhEHGM/GvnVPJ8lYSlp5HW91dENJ5TsjUix985
AMYtHZVY64QqIPRnMHfSavgXAHnWeCQOdBCHUJohLo5sfFfA2MuEfx05PGav3sJs
mFgY7Tt125ggd/1pYdPr0QTH1Ha6Nk746RJV4Qqi0oTiVcoIW347w35VtVrX/0N6
CxCvCzK2t4CC+SUBC11ZUQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
T4CWpcfTtRTLBXnaPdkEDJl3q6vzO8dnBm7W+SDUrYWxsavHCpVaIIWKzM2nMXDV
lpKYqy7NaAyJVbbsOTcjTkKoRLG1AbA1YMKtazMtvGI0TiC7qWZZ/D6sRfxHLPdh
GeuewzUI/bdEyskcf7vP+3kCJl/RQNw+S685T7u1uDQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3728 )
`protect data_block
0IrnDvoHC2smaT7K2eMT6cpdQ2ZnTbNebGkPkUSnfBDgd/mDwRTkNclWfUx8o7qN
zaJjqEoyvqz12LvFqytk4G6IeAoL+ddHMEYL75AC8yFY9Y7PeIa2BHOqWuL42qPO
0J91ZbcBMuY7UURf4eISP13RQi2+BMSL9BbzcUAnXDiuZcKE/hbQ+DsQnM0Xs5My
tIwzkf3rZF3jBuUCFKoOCPMNDWvWe8nVws1BJjvZjMn65GU7Svbr2/Mev27r9A2D
i6S0SgAeB34d/N2YFtWL0kxM0g+++wP/GUofMBv5pdOoGSt/IJ7fqMnFadBpwh0v
PLvy46liyoz86MsEzjw2KmbR62LYRSiJjHStWjJoUKnOExLBeS3ObVadr0WDkV9X
w2ZvW9sCfO9/qlIZxkNxnAWtrWE3nvl0gzOcU+HTMrLC42l0b6s1vH6kFtiKMM1H
hJ1kwjzwVaB3e9ByFta4vef+8fTIq0oX6CYzvDvMJ6jq00TiEZI6OPqdOps1lbs1
Zzv7dZWjKxr4//iXxaurc5tx9QYSNDaImZnpc5TbT4kWpAQQMypqYpNkyuXK4EmJ
Cvpp301mo/2oaSUjMTB0VVOgbocQb7ep3mvJF53sfI4oeeJ4SCC9Il7JFQvZseQ5
uiLnkrN4OowyxPXpvaViuh8HDsvxBkNs7omX1xDwB5mvRza2EB5TYRlEN/CVc/rG
phdQtFI39v4si9rAoDi8oNPyfT6JRJCVJSm75O1cb/Qe9RXMl2FGYIq9hRDd9QWF
pTXGYnKTBuoP0J82Uv2hVpoV0HafiuqII2ExC6dTB7bSxCKg9vDilBky/LLAxPcx
bYm8O+iHOTc2jSuHq3Vokwo5iOWfEOfGSZRg54L1k9597wgXQZN13DNUtWW0vi9f
Qla6euLbLs9XdOhdhoXoaqMIPt2JjX4l+80HuE6I7yDfBhiPX4wcD7PBC4lZWK/9
DcdWTkZkqpZ7qjeJTVBfci0SCxKHOMDjfBSwnHw9F16mYjIBIPo5V33UmNtOwHOP
ZjOGYSyq0lWAdbvgSy5WLYPXlGT2FA/ODu8m+MRvz7xZ3nEiBBVCnj1gvt0NFa18
t8RuRJsHHVBIhha72T+UrWVQjnjTNSSozs2DfAt9kD6x2P4jSNaulgV8WqLTWJHw
izimohHJaFfOelNBKYRzcDGYrYAMFC9cg+jO8sec8YMjCIxNLNp20iUUm2ygZ+zJ
IUp7xgTwpo9pFOGZltET5/3Lf/K/A7a7vv934rAS5w2yaYWnhoDqISU/4OUuvb2i
tUKU92Aq9XfbAj/NfZrTkNcpJ6ZUSmW0M9G1z02uGPbMG5uOilpE4pf/96BunX6V
9SG1MEL1odk/XzvCBXenSEehw//IeUS1r8lBffWTB+jvHXVhVABeNTXOvoQ29TSS
hca6/rIQU53ktjxEk8YJadAi5Xw8vgR5v4wNl4Ob+LzRRCn55O39kZWG2vhUJrrf
Ain7zbbE5q6enTAv81QHYwuZArNIOSC4RJ2tuHR7Zq6VfI7Kj6OnJcGybGka3CXC
sCC2TJCAEH55PbJY85/VlxkfOBDS7Khg9meWprqcM/Xb1Cyh9E30LtExhgtNA1k0
YpFzJniIJJJ2lLpyRg9MwEnl/CshqnbjqYZDXuAyhq/u/iOMemI3+2CMLhqcbUyB
7i/pX77S15WVvcyRv+1p7P44xVyC4qFEQqOXGXJWTj2/T9vW5JZT00UjefzkJ62a
9kVF0gSizfkAJtXOCpMJ5Vky0FmlvgkVQvOus/3/cBnZ99dbhtmzvJLEIWPFnM9z
+UMQ1/sSz8WmzfeX4scQre/1Mfn6dzAlEBTw+kHeIHXeBNAXEMM3/3zXi5BXXvgo
b1BqVlToyA9DBFB6RDW3ug5ZnLdlMyFfCHTfFcJSKXFRzJ0Wu0Unuk/gmNd33by7
zMntC1OF7E3kEgAXP7kxmwMCNXty604bD/YRJ49NIJkabybZ3iIg3Rzr88nxY6dl
zOtLiIrCDiLy9RonyXr/7XgNqGrPA7N00JtbHQv25RJrKF1i0Flaw75QyckrRY/0
qS+MPWeA7StYLnWFaTkMLE4adg7qdT8c5t+rZUoQOJuJcCp45eOC9PXyP9W8UiUg
BwF4MbY2w/EoyCti3vPYwoTg5XliicQUjUbVEodhgD3+89PXH5Fq00gsBkzCK6Kk
Tydob4QrJK4UBPH3H3nV77TNfUMVmKmkrlqpt83w8J1DxBSW9j91csaRqcE2ElBp
dD2OKg38jWKa0hvJVqBMe8juXDPpOo8AqENJ4E+wX41F8Jo3r2gpk3VkQcDJRO19
66lKYV8Ellj3mlBooWR/kjbYEqKIUCseZqSjnPBJoEVJccc3GLOpBIgKfryhWuI2
dtQ0uf/6I7TUXtiXjSMElsx4urHRma9KANWl5e6TwRZmgcdBgtQek5O8yvIaKVPh
tzqaPJIrDphBmJliNfxj+sHXC/ZO2+o9QQLblurYXnGr/q1GKj6WGI+ygdjjkpF9
rb5fYgBKvTWmEpMMi8AJdlufMvR2seQtzerluVADej6uA88aGFBqT0PwdoJNR6r2
Upon1EwwzP7TwTV+enGvbKiKMHOUM+lcUCnc2v7MZitgBC1E3tsDi5zkBcoRrP/R
ihXsjqt/8ZiPT2PX9Ep0Ci3iWpzyYDF+UhqLDzWYvUS5Bx2HW+KI6srBC8E5vCdk
pbVD+9cqcnWvQ68Xb9oFttOv9zMyhRYyJ0MT7hRi4QD5ThUfU2fiNITrJWShwxKb
NpIs2kelbFRK3loSb19ybqkl3Q+D/GLzfm4gZcQqivjnkoCfci3mvFX5EceYdU3j
VbPFleiRW7B2a/3CrvXobRhrUhsujlchWfAHr+bWGoLP2OOPqMXxDxQp5hapYJi6
u9bLMPF6SKbgCH+2fb63XvWh7l1d9zIxJ5XZYxh55g81z9cGDUH/pLT+N2ANLOtF
RMUPDQokOH2/5IOiBO8MjyhTAAXxCTjMLLnMufBAG5CfoUSp/8qOjqX/8tyCI0S4
ORwTH/fdMYTNVaHmO9jmTWoCvq9OuofFBEsSlWycWl5J20Oc5zxvoieTyyqbCmB3
UduJz+VjpgPD8hty/qe2ogcvOYTo+wU6uHYSpIX0gyunXEC1MpUOK20B4Cq+UeSP
x0iDixDtTFeQYwoyFImQF/hd+6l8gnyuGoKCu3gIggH/FIYdKa9sk31FZHH/5NdZ
fTWlFfGtRNeC+XrdpLZB+xF/TylvznH52JQ90WyORyggM1YnE+x1aebn5FAvraHH
T0XpHrZLDdeLYJtBkHKIBwUFD9hTac52qjW20I6jsw1+AXZGw8ecboWMCIHXBKo+
eruz2XxeUvRs6hjxEFR/5wuhC9MtOEiMguN5k65FyCbpMgcoUXqcC2rIFeny532p
JeJiOsDGdfKeWyVEy1tu27Wcq/XiWANL7xr6nhS8/gm8BSmSvh3jLyVvjuTktE7m
c/GKihWbn1Q53HYpcuuwnPg9YJrdI4kNhE1XLDYJXujYw07YO9XbfRaSrcjZ/juL
EwvaFC8p5nzzukBZP35Gklm0ExWpQS11QPxPiGfY0r1gBMvzvsEAxdfSRR9US52I
f9kUG1SidiLeULCH0vCNejSRCeC7lkn67raNUSnl3JObwT5Y9ToTF41VFy33qlhg
GHmLlOWNvUFC7v/J3THCas4l6SBy+UJs5DA27UkWuZHFbMEjnqBDJ81LvSpaxbTL
if4LEKya0Rfamk/haEvmSjuKFVF7XVLxK3zQcRytM1WHq6MKIdX7hqT5skg7JnJB
RjCr///Nw7gIf+nI6RqCOjzEJaaOHvKuKIyRxgYj4kG3P8uHEkEB4vamfxyQzrlj
oDIMkgvmj79qrdg7/pYKDyS1ZwRNFgzf2OEhTOdjoOMW5+hv7VIYIvtUC/KGiEi9
Wi940EPh9aUxk8WSrlhG93j3Pz4Cd79sHH94lws7Fm+z304prNj1fIhz/WDJfJBp
dSPCZQo6u/k8Z+qWF7CsAEvPRRStdZORoVYD4MYYvJ/CSVeeOiJnWFofkXeV9OkH
Lr+5TEoZSoJEW0PlktCUgqBAxfJrfhQ30q8t0BFymYB+hLyuMY/67vAftCvxGErA
zgS1cYrU4Oun9kiU1fAgODEY5ZalHRK2pAADz+NNQlZl9jgEiKJ4bt0A7V6atDsG
KtWCCNFFSHVXdQGHYii7R+7kiL2pFFeUsgrriwMqjk/0H0EBjNyVVOaYsTKxanho
/CuE2R/v1M6WNtFBb/JjobIR7iCAVtOLlUrZsNuZEVpBkdC8DOGrilz05Q/V9xB9
zpe9lrS4v6R/1+0QiSz+XKvmFBqT/M91uAV8xroVL1zfGyFZ6ZGlUDM/WoqPtdXQ
2eBR9XJV3bFZ9/oTwMHURVj/aSdiywrKBAaA6uuinEX97uuYqqbOF/m3x+rwmoZZ
zmNf3vbG19zHX1GiuICq6fO9l537OKb2esXkw3CJBvavpiVT+6Gu7tw1hZiXCa1j
RT2LY9M4Q0r3HO0Tb1xWa2ED/vn4rd4HLucv4oD4PKpiFkLwOS0m7bItpc2uB59a
7E7RxseO0GCySdx1qrJ139CtAj3qBACpTn4qWyUdCxsBTePpiSdWtZ3eq1LjZttQ
xpg6NurOISYyW33N5Zdca/I/G4LPZ5EKWqY90I12TDd9uXQMG0FmY69xbpDVNqVN
f10x8uT56r255DKfIDaUAWGGfHL5pFjjs3mGWBdHqd360VW1+xu9IueratkwBJ2U
eZdbOOG+ds/L00xALWTRMuFjRneKXzG60hB76EQmnkHugrjntb3wtCTuiQsQtgIs
NvgH9x8C763tDAFFgCCCA5SBX9hJ+Z7y24nTj/rbp/v+QhTxwvDwiHejHAEWjMN6
o/y6NLfqaJIen2xM0rHdbhnAcQemqR6gtLmVde7I6ucLaPIUcqdu6vba10YH/JgE
Y5IzNvaz2yWDA0SFfxsm7rsu5n443TjLQYqru0qetHg=
`protect end_protected
