`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
J4tdNBjJb5mURvFE1j4LGerdiYn5gkOFE8RM5Y+fyL7ADqG8DbpHDh95kwTX6Edb
1QjIFG7VZ07Qu7IBZA7iLHx1vPIDMcpAnvPZ9Lq3AjmRBC4v0iJ/c0ZDTMmIphrJ
kNnmEmqCzNTgGkHps0nZylhkhVQzqP7Wng2BMffaZx5KCrJnHoyjRA1O6OSAoo0/
aRGokNPUsZ9Y/1EaR78fIQrNFC9/tQwjSbOa3Lq2Z3Y93mmqkNkjgtZENUCbL2Ky
7lgg/0ReZUrgzNPBhyh31pmFKNeYEvUHv0Wv4fpVYo/05XMF80FPi2uVA8vK9AQ3
6jot+I6aUHgJ1rG+LidaZA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Ax44dQZvT0hc7/1tS32aYidgHasm4+Yx9P9mwAslZRZ9tgnHNdtGyKMWmxYu+yat
L9aHLl9GUvVSfTkbw0tw/mHjGvt4VO/01liFkHF/jZvITLIim84JumnxImQBp38P
HUR7saQvXQQ6EiKQK93+E55z3H+L0aTVyQbHc41uSpk=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 76912 )
`protect data_block
vYSBSoD+ZU7K0Qd74vRD+DvxsD6sKz1lkSGnGoiMnxd53RnMg49bhu/NMjkC4AM9
d2xO1PEcOdBsJZST3sBbHUhdvsKVXfowPppkx1QQRrGjdtR3i+NgKizs0jKUOxbR
Ev0tiVRgYHGdzTkNpWoi6bOVVHPscmCy7mHTk3qFI/rG27quZ7PY0qFwAt+ONZHb
WkpNFGjuSMT2NZMwUobELcyLAkyOWm9u8FMLCzXnXDnP/o5QPb4yJJFCKwlGTqEZ
D6RU+lvlm1gFVHbbnbMcDte3PVZgz66NMiBr8ULHlPO9qJpUrnH0R8mw0Upf2RCI
2dwS/SvhFnPoboqAs53clXxDkFLvIywv6wfDuJh9Sw3jMokp4hRmEaYX8LkBvI0w
JzNtZoc2GywVAB8R4F73D2wSl/jxgZPQLXqO/WZs8i51YPGtFOhqdjkJjgRHS9we
UiopYYwERyN0mKElj5efMXG3Il+Y+qVq693TBa2GM3XMLsOLoIODBdI4p5D4lOoL
nGSNlSM4+4FTCWTbzlFNB0cYuphNRRNVj8iq5grymx0HRGRl3wdk05zVAfsg6xGi
+t6O4BX2/SkNSXRShP9ZA+cPCElccNgiBELTgtu5r4BGRWS1GUddRGrfB7brvN8l
hT9bSmiFL0p7hYrs7DPglpi64IA6PUfW52CzXiqlW3MmvZAxupPTdFADMwHbiZnK
e6LvbrbjWJb290SLI7tQjIKsHmuJZpaGvW+uQytF2fJGHUCryUQa+UGtnk0dVomd
lYChMmCfFlnagCV+QT1PtqeYPHXTHA1yPfQd9IlO17vQu9AOTMrY8wjciOarlrBG
Ao0PL9QZZVzdyV2fAjzaFKbeGLQ25wf8NACSfNEd5B8wI4BpvJBde8Rd2FZbwaEi
cOm725du7iXbKL1yt08eefEAmbwVmwdsrvAQnSWMCreRUhiHfn3ldKDCHmvZTOly
aDZI+1NlvLtcQiMHyN3YBPslW56RfYYOTphuSZejltAs8xpDZx45NTptXG1lBLdd
OJ5r9n0AlEIXhYGPvgJEAH1Wbyp9ZDM7SB7NIQewyAY9veF6nBnb8hjm7NH/zxCO
6IAhkB4hFVrBOhLUfxREOCS0L3LTLr8UOcuUWWQR6Aob5YE4CxARe86Xt7jDccap
LaIWriHJ3dU5ykaowO/5sL9XB5ZpEYxrVEXEnfgHfNpxyevK8ASpSzQdxMtSIS/1
tkfhIuyQBWQATXbPuR4tKTPz3J/CcJCdXGLvse2vAuN1LyjcnOq51mJr/JpVDPaL
SHnw/LDNh+tFTYq2J2ZyUxOub08jVFM2MVVWawnZBe5IbnNKO0CT+dPvdtDJbjCt
waItk+0LQv2bfxerkGE6+fXm8xRJ6cKY6glHH/rj6rKbgXmvb5coADwNRGV6Uz6o
S+D4gr6h9b2+q9WTidl5wnGzb449ijavIPp0L2dhDZp4w4YhbSAeh0/nIDepANBq
Zv9fimaXEaFJB6T1rBLE90KelvfSNAok8RBOS5/VosB3Q0B2pP/0fRJUqIPHangn
KPh3H8SArS4hROKCmdX2yYgqfb2lz3Lx13crWBLT8PTFsxprm6HGOKPH+8KXXDCl
82809jIZGBHKgTKsjr30xZg2Ij7Vu0fdtV2jH6+npB3YYNSADhNct9NwZSxvm5PK
197BuUg1t3LXu1SRmnVjXjCo4edE607ZB34MlFl2Ro9anXcI72X04JsRbdtYes7s
y9IPidrGKK2I5kaaj4xBjBxrFMl+/hIFkZ3kEbNp+yCCWFGrK8vWeva7Loyllnju
PLKu4mZKpgyKkVDrt6UMdhGatgHCcChWqPDn4+hjPL9RM36IBVjE14ciByQAg5vO
/Xp9fX6BQ7d/a1JmAaiRkw5eHmX3Liz8OtiCfjvyEMbEYa3w7JSjxU95CO2V0cgH
9SvBo6tvGBfi6tSbTEpqIaSLFAHdOJS8jkL32DDc0DZ4rMCOZ2hiLcPOaROamJrm
OfCjjz1OZokdcRdk6YkrOsInxOjFIjMm3DHjkihEk5hRLodgaWxcN2vtMm95jYN/
4tY3xoumzkMG9wvinDB9HZCM0aJJ38dem7eaTOPGqohMx7HWVYbR2cRgb+ZGUiTP
NhSGzQ4m4ysQwVoQFTf7vcAucN7ciwfkLch2+Em/8s1IWfHcnFxpAGT2zr6M09QZ
rucUDoEYRytI2pdDmsLLsQ6C7gEgF9htszoRo+ApmPYmDzQdt/9Q+wAT1M7P0j6X
qn13KEo9s7Y4OSPy3WuHLNq6yW3HiJ7QUq0RfvWewX+or03ZSyLYi3JX4Va3U28P
fS+mnR2PEORUmb6ETkpILRf5mebbJR35+A/RjR3kUxtttgiu2W8tcayZ+Z9JKSgd
qOHuZJgi0H+gWBaiAOFodMwubUAGuDqdvQxxJpkZi/hQz4AY7wu9R1ff/NBtFprK
OJrShSLhnqwt3C978X9B7/h7Y9v7tCI9vi+Zd/VOcC/Q59BiikG3iJPMMseLAOu7
f3k3DJHtakt7+WOyNfUoV5PNPcBvlbRfwnXOHYdihZ7mNoVHdSLqXYVLs23jzpOz
Tx1uJS2j0yQA47ts/1AtaJ3NzHEv7AtqpANr+l8a1O5C63vvXEk5XjQA6lhcUnhm
uEk6vrtlNPu3+BsckkVX11UPqUtLZpm6/kNF9STliciLniy5K1dfs2jSOJ+aIG0I
0ebrDpriYljAXMm0vwhQug85mM1ltqHp0opCnaop2d92NAiuHW7HU3xlhWqgFubG
VQcj+2XUyWiMqlQNSu/mOUX1+79UF5HeKzOHpM1urJSmP4SIs46NgaigI/XmEARJ
xh5+MSTGArO73jUiQ1q6Q9aslnibMbuchbyLix2Qnyx3ZVkHAmZi5fjqPaMKkMT8
jRtP02mNawwstnTelZrvGzV5ln8H/gDgEypGqtR+pwaOGsq/an12VpfvFnfJMCXI
3ZsNwLFedzLJ7wVPivv4HmKoW9UYt/F7LvokOG/asFk0eojJCsiwpdq3LXPyDPfY
M6391zHONncShUu6kxtNJ7je8451R8Az8AqQ+YcvmslQksPWKOTrpFHcn+HYIxW0
dWnxyFB+TLY9Zj95KnxJ997Vwc2yD3lZybzfRoA2RyawNzugNkHh/aRqdtOk5hwh
gSxKh692417tPLaZxFc2j7vGMpHWqCjoPrRa2i9Wjb+wkK0hX/cFO9wo+J3/6O4r
783jP8oCCzu7luNf//k8Gt/t39m3hjXSs7V+klV3qPy+uE47Kotzutv7iZ1zyHF9
lID83inOgsU2g4qbHCKpNAskUs4jIxtJkFx5mmjGsN+mu64DZgGJZj80DU1H3hl8
a7Jk07EzDnzL6NXWZcPtX4XcTTvTgL8/oEaizhPsz9zTJhC1Kj4te2dOEZ9nXeWb
z9bvgi5J681LQvkpZxfa5THUdizjzFuL7u4DyF73VGjblxVpRvBQTZWlblrPzMIS
vMobHD2c2xVFOwvBgfScdxbqIj7A0xdl8a0HlJPa2UeSyeSc44hcJKdZVuupdYgv
HKpBJX9m5ioXMGHsT4BRRB3yFSVoL2hNCUQmv7ZOSg5d4HRJwpoaXqfPO+qauIU5
GXnEUMAxgcmAaLvtvTWztU83YxIOGpwr9MNxeJzJdfRN+zn0/ZKGUC+aVoSfehCy
9rXw7h+raRR5RVLBIdy4CE5rEaL2+S27hnwvLttO5YAxn8pB90frJ0YRjR4XxTwy
FKRZbyEvRQqmzE2xfDP/cGBQxRCj2cypYblnP0ZQry//l294Io+6fTABwrqasRAp
rv7LTizedaQJwYfnG0Usg56LabvMfClNp4IGWTIhCQj1euHPrBxzyQxlKY/ezJAQ
IwASlcFPHDu4IdorNiW+gkemVG2dyZ5tgrYO/JZogaTbyjutUgJo7IXZObbPxtBy
F9Sujkp9CVIIgvwXLTzvFZYwqEIDShoQQXr94cZHt+U/3oczh++wGMCA2QWgwSZ3
x/0AENRKmiawQqGNF/3nJx0arlZCUJAq4ERcKNlpdBYygxtlgMQxZ/tpVoeRKyt1
NNg6N+QXLrnCPk2Z1EkLdHoDjVmOGzSwj28WLP+On+sBqljNKSRbN3iETIhdB8AY
ViJzRqT4ZDW5z/IYEIF3ur2RHitOzJ2aXmnmmngDxbfKa5VAP/6BG7DugYRoBsp6
Kj2yTcsvw0F2aosOwtaY0SUk1Iem9kxN4d4UjQjnoy+DL7rj0mCCb69ACtfnLHhO
Rg9Gsn1uvpWsulmieJzFfgD4bnenEIF3IqlqshjQ6xDZwAQl/mqh12aCfJfuwraG
i/xA4TY8rC0vRTzY9ttlptt26wo4ixqxH1GAjwLA31nwm2RzEdlEMZ7Ysck5dXYX
JPrpkHatEW/Pb4BDQfAkUFwMjowjyT7Uqhk7oNVwVP5FW3BVax/MX0ynyH9jENz8
PXam2ltucqf74blLOB9EPSV76JXpR80u9b/KR81Fl+fd8xw4h2SsbUFrH9s7+qUi
j506DfkOomBsGhWBLkARwoUoiRLKwbkxySDeCTCzmj4/oRlkpJXCDYNFoRZVrEzU
5PbXF6wNU8YW5flLaCWHtXTSGNzu1J0uL5iWmofS4tQBBibdUtESFe+0YctlQKQ2
pusjLyf9/Jt8tNUQxzIoZNUYWTAfErHYy+rdxc+5plTTA64TFKfa8Gib4r1CohhO
KTjadqaxC0upIsZVSLNqPB8mnZzk8tGm6SHw1LgVwK9vav3ELecq5LjbpGQ5J7Tk
U0ge2Q3cS6kcQvABGfIdCFWvDkMZjaPr4znbZzMnaMTlLFFKAXTp/fpEcdEOllWe
f0yaPjILryrhE7uAgLHqenOK5X7XVo8fKRMBKzGRilGFkeVPw4pSn6Fjs1pXcTZw
yMiiFdX3eAwnF5aiGr6Eu0ZKNn5sxn1lq2RPz9jE28qHFSx5xbl94TtmfdE+7E+x
ECrHJaLvqiVSQ2DGXaVu6/nxLFTnmiOrRmx3t38hNv5x/vunyapF9oMBNpVzobfF
LIBLZw6ix1hC94O5w1i2bJSJhaS85IiVUIQ45vCeCt8ju/2Pya1ZsOwSLBZpcC/u
vRqif1hk2djN17RppBlbmhy1NVw/gktkhZ1HEiEdeozscMabSvpV4knZI0pz04lm
TyaEg5iIUqcaGpTSsPDL6Jw3zt495+K4v02cvtUITCbgGvLmjoyjTLm5Z7H6ERmX
LGPuRNifp7p+W48QzwExnbbHa2FkzrAf7r7fWOwBcSzpP5fk+sjkcHU/OUvPKGkc
35/oxfadjUjLVE8muJbxZUCE5twdfp3zIVGH9It8fnABByxltXMtyVSoK6sAoQtT
IBS0QXCFFEpmpq54KuiU1luDyn8mySXLFHkIwrigwVfhh3JJn53qfwy2fl9bgEc0
IAo61v6m0pdru7oOi2utCyZmGVmFxYCd1t56EbiuYd56rRvbrkALwbnORmvhWJN0
LNj/ATh12jf7QmIHhwDHjwwTQJ9FnJ2ykV2dwBf2flqEkI4jl3qNqauTGtb3dyNh
o5WW/r6Z0QkmZuA97w5XKto1S73Qwy7dRpY1sXw0XOhYYrmGCKXEeU8sb9WGMSNN
YOsmcC5elWcdo7xXUBznkhH7VoQLasBRgMmbqXToCw/PW0uH3iujVlSHXevMLmNq
6wMOOoLXbS0RCxpf9B3BDjNiGKQY1xwr+lGEvwL3M1wDbW7gKo/Vm2RGdQI8hEJO
78cUBR8BXTI7bOWxR5JfoCDGyWKPA0HvKTiQoz3BzGDp3ADP3ve8PdATaHcd6NnI
yiMfREP5grcqemFZrFCvr0gRBIynLyY/rxaGU+RTpIJ1Z5nr8GwzGOjAN6h7iNkm
X7LLk2NtDTBJsrLFM+HaEv0dPHr23MPWPANVjSwAyrNfk7XtTeJUeUXb983z36eC
h94PLYVJF7OGiybGaJ7MIhIF90HVJWEw5NKBGBGTo3pSXnLhc030N2B28iVFystZ
eCAjxYnNfU9Qv47Gu+ZSPh0t5Nk9nJSCqqFOFDz3e7aRnPkrVSfQXWKeHeN2Uc+f
e4ZyuT4y8tvrV8zr0iAAuY0LpHVMG7Cr/snynvtAIcaCFlU/FmYHTpvZJTU3ftyX
tZE6Le8SPlu+4ko+oClRd7dBL9b2VlblATM6byokga6ij9Vx9pptPD47H09hbJLN
1b2ykV6erLEFYGLwegGvFQbVZ1maUblZM8D/8xVk47K3oiHgY0YHXannBJF/J5VU
soAj7WccCiDQHzyL25TDGtHYrsJEfYH/y872dXCZrRaYJUkr7Bn7vZSxp12xfNjF
iXt46GKb7r/CHQ8LO3fUkF/1mwRjqcY61Gl6OcgrBB8VthNJI7iM5zBIwT3LMjCu
L9uu9QnFn+kSwBMOlCMwRr2/q0dKnOM10ajsyicNXwYoLQXfIhjNXkYtl+XRbGAR
RSkLE2RUzj84T+AUigrsmnrdOlvew/YPRBOg9c1WmSaKfHoES+MZ0ZkxKSdzTffz
63YAPr5L+DUdDN2waNJSt/aJ1aVeJ5KzpSIkZDdmFUN4+hdnghhKhNKQc7k/ecVQ
yTEJW20pPyQ29eP4lattg2XTbj6Z2EfUgQuQHTHrh0ZdaZHUnOKHEIJK6i4K8W3t
BVe5LIFZuU8xnoY8QNSFjJ2+spHcm0ETRmE2RWnWaQ+gdJOr0fm2rW4O+rRrDoim
jk5X4jV9OzZ2h4C3yEJz7tSiPAy/pS+ibaY9itCINrzCbhDAO87IhmdXw/45dyPy
jZ0HYEpU0hessMlZWZSgpRxwzD8Il7WrmxhZkOfPgwuX83f5dv3OzfR70trXnPE3
GlDztHzjfG05/iQ8bqwkqKs0qj0f+/bJ8YI/pvkGLgdliz9x48rdwNsHX9bsmCCp
Z/Zmc7EUaBtKh3zULWJi9dFw6IysnQcEQbz4f+s2O+11k/RQRpMpcI0O3ygYKK2d
QbB1TmCkxkiZwJWjveYE2h0RIC63iRCCqOOnIfo7+vsSRkHNtQhBMXDipuHNatfn
nIxK9f0aFW237nocqVKx2QNm84ii0KnDiHMyFlZ/XjkZ4Tl30yjggQDp8Db55KHc
8QIHzAGiKXc9JFW2jyQ/oBmxagt7a/vKrBz6aQSI8gyYB1grVa0r4eRBnrhAtSVb
RxCilZwRZdYssBp3QCatJNu0sISoNWXvwoJUdu2s17n/ng7A6tOuY0Z73dsbqB9+
TrwryDcawzKogATH/hmv0rsxAzSuen6iPBg7jpupWwR3eKU+gyUlJFxFrXboYMyw
8ye4StMyaOdEC+I0JR8PC1sjHALiohYKHC9zzQmIxdhSYJ9lqYvN4j7x2lClyz63
uoLJ7ccgMO4xrak8/cs2tGCY+yD9HKqkSngkYvMQpixNm70MZcYEsGQieLq6Fn93
kXb+M2bxZxzmZUB03yBdGVJm1AVmwn66YGBEXDPE/C0OEWvi2iJnbddTNcsnSkY/
oDxoTipb7PCZgZl7FoMcKXTwA0DVK8PnjS8/a5tzUMG836wofmfla98BxKg8rhh0
m16qB34DY8ryr2Q0n7tLdkE3hV4DhjwmG0dwU56m2QbR6ca67WEnyXktoyG+l8lD
3J4g1DiKFQpMONvTN1Vpnpy8qHgtJ+f1uOUCk8J8psKp96Bavl79e75ZpIs1k4vu
PWQD7rlDnhaJLfIuHecKL4oqkiJM8sgGyonZdsvQLTPTQT1D52aIEDWCEHXWoU7O
Ol86TaWQyqvvhPpyz6lICXpxh6FGhKIzZsUcN2CJpPuqQDs8++kGsfVEO2RQTFYs
LwS75qTThskbFZ8+2Mx6wIdogLkgakix07cx5jdX/0EoxsZoWuN0DpMkOYRS4lks
YXBKgy+n2T4I/0/q390TDocoVZCCCW+QXVmZXJec6FvEkjErXatVEHNNZP2vRpqT
gneL5K4XlxnImf8MT3Ocw65sRp9mIlEFfMSuPIFIV3iB2XH5kQvPchQeZFLX58uf
aA/gzuPUTbCSeSgvXMv9jQ5Js0zG/vjFhHdNDXbc+tR7HSGPGjAhSO3y5We8SMwa
O9m4qhHWhEEDgn/YNvg9QqPyaKksxseIEzmOhROPmcMJzrh3ZOgeqmSlfhMmpCPc
p8BkuIyqaKqv1FXUZeHA53YBREH9DEfC/Q81Ypwcn5o7T6GwfTEEwT/Ctd8YUDFS
LyPwvrZtzoTnkDGOoVZjREPz+jMGKixgxMFUXSAlclIl8tVuEPfOJNO+Xk4wP7YL
0KeIsyZismLKXTuBleyRqZqmqIGMluBw/UcTzVYA/u5IyC60VVQIPdoTDgWwg+HW
If4ceP4kTMjqc2BuLmnLmifYzsoWdHklx9BOj77m3HEB4f+gpE6UEujXcXZVhbFd
oOzJT3+dSx4D790U2KXtRgxK6UX7rXeAbDjyh/LFoI41j9MrbLGx5to1g6GiNTHh
D89SaL1i3JnZzorcntRgyziNPJ9atqIwBO6mbQ+JNycPWsVR98rvhvsR7JUFQ04P
ZndcIrvq4butEKun7wv0xiTyHrZ83ex5cixmCP5uBEWsBpNkchCKN+xK2b/aMokj
cmG/gkDH3xJhh/B0R4Ka/mzzxY+B60/JYILTWXUiQCxztecAWkQCiCG1UIv5Y64j
uW3t0uP1+PI2JaB2f4/gDnVdtwzQ6TqRVnF1uhvKvyVs3zXNcK7XUzAMT5qdxLHJ
/UmFUbkGkTCTScav19YNU0oBY2i6w4Aj7FSpC+17R+1Hg8uiCPkZc6l0iCMwKW0L
BeUuwdqcFOzpWVyP/OEFTT/UUBEQAtI3apl3qOMg3cWpu1LVaLYGdMkHavcxoQp3
EFoPiZ9uKCURuuccDGCVm2/yj2mtSUnTkyQnPIgWEv7H1WahgQ0DPxHwsKq3Dx5a
0Yedt8/mSJqW8RGOfgcGhjPRKV/eA2wnT+jttpVlcM67tEv4vTzQEPVhki2pCjfk
SQpWof03q2D/g3r+LnS8586NflILw72CO+crDPfEC+au9gtDJl5O4XfSYuf8gbee
N+8v0jamvin5P5Fl4jRBds3h9Nq60A8WjseK2bjdGwZmUKNT1hJ6nZYoDH9vP7I9
7bNT9e+4f84uHVG2EpC2ZfzlvlCSdeY9cbILKDiMpAYBVs9eZEJQfSk/qsAWIr8C
9fXOT2pdAb7oPRQl4KrvOKdvMJN3icmio/yNYEKyzvE479HZtbt/jntwuvwUCjP7
q5EJst8zZ9yJVQ6kWboc9hKesezJAaXXqZS5pRbj5fyRxQ9pP9V6FfvLEGh5AvvZ
z3Yalb02DXPcSpeSJT7dHD8D4DFQJKdD4UihYDibh8eOHrJz6zph9Kf5DZ2FRj3G
lXuSgUNRl9H3TfcjmtilkgLktubkssasD6AwjXY5kv3z9038a7dLp9f8X4k01zcG
dxCKQDDdNgE0kL12JX2Pg1uBOi6O8wj+FWBv+7+8YC7zZUU+xPQl0DXM3iCnKTAE
3F4gzIkMyK4jbXhg74oDSolnIrSpdU/dNFA3Fdx5490P9eS+kwCq8Dt27IWgfcaM
LBTB54v+ZWh9D61nNGCqg7A4ECxsz+jzcx5/dtsY3QXDAb+9PHABW5NxclF/rfJa
v2EF54mA/DvZjzVNkECNum8WAAQWGU7MoZKWpvP5H7r7oAaoiO+ALBMP6vlEqXon
KG9bxlrntKD947+JLvtod6Srv1UfQ4/USPvgAw+E1ICzPQsL5aZz2BbKm8nnBlbH
tjrvQbzKbVQUVfdkdtdppGb+J50aFCMi6Nc1QkdWmm8v8iMqss3BB9yhKofYX8TV
uWVrI7rLVpW7fAdt2pOCma+tKsOye7gCdKdMJEsKrGvrOLYkgkAj60CBi4t9JBNo
0MOXIW0+mGCXp7Xi0ENZ6JIoYZTNgoQdaJK6SlW2DYBagq7YrwbTUO4oxd5nt+rW
ahBtgEPJwnikIxnEdBACVy+YPLWqsas0iQSas0SgUE2RGXM207bG/UjRyCS+8rgc
EwNRRV8QI6h+Btv+5mi3DvtZ7qfNSvlNvaQn6pMEThdUaU/xoj0JkOm93K1m0jNf
n3U6VHSCzRZTL0QqAy2YpfCQYaVqMqDhlqJHYKnwLZ3vh15JyGkFBNx0OEZqv7EO
SENxgErVsW6lWAZwl0oiZT2QlFJUO5ZUTC/ToYseXpfwrVgiW2LWpIlD/kLGeSrh
isRHqxnbSSNkaCv6gx0mlzXPyAVq2Bj2mz/76Cx8NPu0MSTijsFo1zBxEcYC36lw
hgXr7KqBo1yhL3c4TXaQsFtYeFyjlw3gRD6leM1rQkd4bBuQCmuQ8b69gltv1xs5
Ps5yQrq7Pk1+p4L2Ptk9PprNCCTgKEVp3drPi3q6e9YpLlKrTyLmA0CEYqlVt9ze
odLvK57UKKtIP4B+Zsx9403v+FdE/fF81PkXc14PvpF8m+xUWdgwAYw5CS6VAXRG
mf36R28JFwnCsJ8V9WEo+Syr2lBSRs8PD6Rc50kh/6e6CGUOc0DcPPH4rvp9xf/Z
pj8FZiwAReVOTlhdvvibXenAzBZ67kFmkVTilTe/n2109m61oiRRWKp7e3nC/QRA
PE+OWBBGXSF2YsqMWQ6zDRmhQiFbDtQaSg3mDd0lEZcFvCdfYEJqTcWfY4/NZuqy
auXOP+dhZ7dNx+P1k90ytwJ/SCLIG/f2iw3t1UouNcBK0aAKsf0iBQ2SL5IMdx6t
mZb4zbopLlX8X1oN8kuZULNrlny/bcXULo0m78nnCi1yIlK+yFnFWhemhAChiE9R
hI3HsxIBs0Q578dyHdm0Sm1L0ynkPLV+EuiAvpSxJ74Ir9vkTjT7+Cxbr6t6bi4o
ZrwjT8JXOoQQdDGeLE114oprCd3MhfqXU303Vqw/G36FPs4O/+CsaLiThDGpgR4A
ylqVfKXzJBmVh0FyPb7IMxK7HJqYfPVGR8ripihJ5ayw1JFtDM7j+0j1WmRs+hnn
M2wMz0KvhXwclJzL6LvJGyBLhb6nlAVuLyFZTK9ZWh+S91QHk2FyAk5oc8dmI/AN
zfTgoeV2OBnSywVWW+L9ihKkDD/Ul1lBPumqIQve8IZOY3C7XPDqGcL+K2pLEp0W
wsgjDOsp5IB9Oy40Pyb6oS7hbVqGA4eYeRWbLai8cG9IDcmok7FTTaEmO7JVP4KC
zA3UeU/RwIo3egOS4Yy8gbcv6cbF2WD1qT6tzZRjeN2e+9Q0E3HB6QrZhU3YKoEZ
GwV3i2mYW7+WIZcoCucJZZIt4j8t1bRizSja8gIq1ojmub62p8AXEHDxiVPj7ruL
ATu4/GEWTmmrZ829gB7dJoGTjeFZqQYrV1zkloU675M48+Ok84MAsp/BAroNtA+3
wnFK6iS8i7Yu4vhvQvTeH/Opg27PZxOqHt0dSZZroOcUKq+U4d+2hi4x0Lbv4ETb
v10GXZtdstAyM6TL5habA9n5TTxV8WzbSWj9mnHMPy2U/oyXgP4GjYTUC/sO+EFs
J899SieJtbF6gdc6OIAgX5qoTeB5v3HafViY4Rnyl3r7/aMcSqaZOQhgcczdCoWY
k6qi6zcRoHgP72ezh/NnCJnkJQJnyvs2hQtm2SHlsaO3he9UtWW2OEh5esRhpDmC
b9nCTT0+EfA+YbylFD5QQhiWI1Sz338wDFXzp745VrgL4yIMFt9Gukw/+xFqePuB
qKC3VDvhHsrkGbGTKEtSTRfLsdaGZjRgEwnadN9ya+SHlZ8h1+garCqat3Tl4erY
G28FTNnMVKXOjgDSZ5E8ane6bEYmrY+0L73FoJLCu8iy2e7mdRidAmTuZ22w203P
4FqzmF4P3PcAwi3isEIhQIIxpKZseYNDcKfdtNP6H2buu6CwA8/XW9Moz4owy+0i
SKFRENaodeLbPHK4OIxCcWiLZL0DuAOD/08axJ16CL4ZOZkvD7G7xZdGnwkx92Je
gUFuzeL6HTrlst52sL0xfhABskTuZXqk0GomXOGIJpQqp2Z04WwsDMXe6odeUEU/
LGIBB5IbH3YkjhrTrwgXAlr/ifGu09VZjh74wKRZEvzoUT3oEW7D/syPZdfylkKc
iuYpJCK6Cjy05d+ze52PsLugYntkTU4C21k+uj/VdQmBaSefO/La5k9RN3WsdxHh
uEse+UNhOzCN84re8lXsVzSVcLpSJa26/usobuRHlICQtJibaHl+bhlBKsVh9PIk
IXziwM7HGTBLy8eXr/GZqOypdaNY7y6Jqm7lhmy831E1F7fNtmzk0Poe03aE9XEf
86WZDBBndEOkchtWl0TEEMxxmlvbhwGidxXT64+xTOEwKI1c+q+GTllvgXUfODgn
v9HQEW4TglIAMdrH3bjZ2iPoCHzPn4Eq8Wbb/DoXbSFUreuw6bBYPW/ap8+spLRi
dSoyz0mV+0r7c1YjoVQTUjPB+ZN1MbSX1870H8amOJX11kbBqjuxl3Xyb8/TBCH0
mfVut2H2mtlxyKKQ/p5cz+DXSKAlfFx7D2f7nx/bgzxJetOY3KWUi3GuuP/qNH6A
AB5jks8PgfDYR9q6e5cxvhCgv9WFsku9itIu4FoocQoCnWmewi2hsJJ/HmFbBvaB
blFDqrw4V7Gmd+eyStiv74PBFCvlHlylWCSrv2mokY2xU0DxhozJJwy6A/jISmYY
GEX5wyGbNFSKT2kP7Byn40ILeOr0sr/1zPy0En8S8zMUZq1CbpLxCHtIopGUKFOW
6XNwjkisEseTB3qH9i8COyfaTE7yEfPAHwouoTL06rWZhH8xvj9cLTvGiVSjG+Q5
mVPN187LWEGkNQmC7X0+akqP7927F2IOwd4Q+Mxb6EU5WwHBg1JwSggpXPqPzFIm
sIkfc/1J8aCrN6t1WoPT3V5O8D9VcwP+bEMH5giW85HllPH77OgAGipt/Plb+QIn
OPLzYW6tplpFD+7aLoKbO5KiOP5VsjooVtSwf8/X56vKwYNoB6Zw7u/uXkQ+aVhb
p7KVATOISNwuT5O13gEbf72mn1EdRrxrKEtmQzadmNa0tCIOs+Z04vZMG3aP0BZL
QPUejjtnLyUSDCMaHqk/6o2aFHm5+C3e7F3FtdL1OhJpqC+a4E8wTywjtdbCV2nd
wEywn/hakycvdNjqJr09jo/bkSROq9mHaML9cep3SvHUkxtFYzpuz/vsQ9InbE7F
fh4t89PAI5EA5blpuEdmO/x9VCciWC97AqjVrwraoWLSL6USqmVDfvnB5PnWd5Aa
pt35LtlhieZ4+1D5gXTKCbkLYRIg1jVPyT6PAnpaIodGyF3xpsn9nFwgmtEK1wfI
U/2Xel1RAgJjv18cQqAu4IM0csE5yIsqYDTdOexHTInQX9s86vKKZf/ZuXRddHtW
MsoqQUC+tIDpY6o/jCk9YzaIH0vGpP0EeN7jMKzfimJTfs58kacexIWgCNDDZoAX
5q+SzxeFmmbVrCPtl21QCmLr0Me2/f2MJ7re7NfViiXNSw89f1NzGeIm5Nmm4m4u
JVBx0Lwuw9DvftiymeWGgl5HPfAe4wkwoMuFZ9WlN7/CLIDFazu4iz7HdpAPE9t9
buAMqXeRglIVimi0JY1YHskVLAoTSPZQWVCANNbTUmf0nUm8qRx/EGaGy9fGE3b9
cyjDs1gckIMocedEQ78c8Fc/XA9r1htUkBomOEk+XQAJi465nq9PHCm5BIkWx3OV
mzWR1hZisYm8/H9O2xYbHgrh8FPY4YXPj9ogXQATvlvDOWspK9o9ijyOo1teexjK
67PiG+GYJ+/Al5oAd+URfxo/rk3G20nKzmZTkQTFtsIJ2S4a8Zoa91C6EP6mqegt
l3GS6yaZHiQ8CpIDFONCLWrUMId1RVlaGOkuhy8hJpBAvuMrz40HLxH1bbGu2r3N
S1Yh+rTB9/sfcqLot5PfD9Tt+J93cT7ejdDcn0DqOqC1ddwD2rQ5FfC9rHch621i
xGgrG5kI+H8NlaF59edOVM89vijgQBRGeTGNwZcx64z716Ghd3gEuvkTVf8ueQEH
Mh8A9XpjCDFfh2UanrFcR2IBM1Yn0R7+WMes5bHaAh/Nf3L0pyaPw9k3A/H489Mm
ruvefk3+4PgkPfgeJE23eBMBC2PXDVHaHSV+ypWflpOyU6q+G08NHCoAQ5lXHkP3
B7L0JHuvi3Ip8hWiinNgPcOxt4ch50DJ9xr5mriuoFq8MYFXFJZzEIMZQED1hZ45
PogGvyoJG9LwlRtWoEbH1DoaBKmPM9J6pIE0rGX4WYSA8Unx/N45W9e3iY+/myxS
5SbDDNWnWm624JsQatL2MOvuVZ0BfbqnaP+c0YD3F+6Xb8nUCcRYCZT6jy16JjJb
ut68RHivkyDRTDSswMgTHM2a8X25Rl6fsAV1a/rlVdR86wPdGFb8CiadUaX2YLxP
kPzU3FyoDRQHSOeIuvTpvflysrTaDEym37uBZBnNwGPCLiP2xZTR4KgHjwHxIbqG
yd2D8BSLBFfF4ubP/EjChv0pAPQ/A8n4ubAvgCzCzysCroN6pT77auKDdtmgkFw0
FE6/LpTUsMlsQOJuZNhSsH7qTQwxGwMudc4DxGEU5til26g8yVx1RYOiZBJgACjw
fiIyLpwN1mwD6y3HXHwA/OMsIdVZ99ddIIqkM89Dfo5ebGsKKGAg6aYaIJFS24Sl
ObMK6Ex5JQbVAmtIkiiiJ21OlrUozylFQkxHxvWvxzcrBu/kwczopIvDO/NDyKnr
obhmE9I/AfshSSY/FRdNE8pDlj+DQPAJLTiQu4aaCuAaZz3M8d3rzuQ7NG8uzCYV
J6cELXBZziyRvGNqG2Uv8oB9HMXiPQRqlKB02awyYe+Q0nKPCrJYWZavpjKZGROC
3U+PUa0a2kiXkNRdGRjotdVZbI7C+yuLGuf0pVJylPziPyM3ZNU1fBtTq5Ap2pGK
DESdE55gPc6Mld5zjmiQ0e/3W30AhG+ooxzf0qtGzDIBP6WelX/hSQNXMy9eU4e4
CGFTdd5iqsEYQ4YYmAlrIuWSZTsC2kn8DNC2T5iKNxDh2e5P4ea7XIxqbET6hCK0
SohwrI1/r2GVVHZhsf0l0jVGdOjgjlU2zuZhfphCJj8UM0WsJALemgoAXZJJy6sB
o5jlDERczeo97QGGxqOaTi2YfUHQDuIHbeCM+AZ5Lyb6zvNeRNwEYRKDRgyXXWcB
CAxMunRI3yxUFIurnHiKjQz9MTr7JLJlHL1NGYJjqWHs2J33GXfvNupuO/IUy1PG
ONj8wsic5sGV2p7um2zU0CXcCVO2vEldQfJdlVeJN7+M0S5irQxttzmfq9wOSueg
2qR84qwMpeFL/7w3sNhV4zahUkpfAg4I+K1KWtEIOGu+bV301O3CwE+HzlchuwSX
hM2GNbEgJp2flq1cjKXK/VPL97B6BooTi50yCytXaTy4tC4NUZ268ILDnbXT7ATh
YA6Ypr3eBcJu30KfjYcmGFtAvDtOrh/V9qnt+YekvUEyfmu8qLUYj2jFBHTRvoD9
j0uqqRzlp2hEOjkwSYSsQYzewcv7v0raGt8MXHyl/4ivGnYXsZiN+DGQHJjlnvO9
oxS1n1eBPxB71KYt2V7VXwyPyyp0UfYDbcUIcm8MExi1N3wTdAKSeZ8VL5lwnV71
NGul+ig2MWWU7QXf/LizYvEf8fXOWmh8b0QlhgoM5cURF9FmPD2594MPPZtkl4lO
Xy2Ysj+RIeybJ2+BwA3i1yW0mj5tl2a9XA8ipw5/BdXxTtGXjEaRC6sSSzsw8tQG
mQCXsFtE5UBz0TH3TJgE/8GqF2vccOSBDJneDp142fuSXgb1Ivn5ZcQpByjCXuDk
FEu3eGpz/jAGVkT1/evYwbJ90f0u2CsLfRRg4vlfVlGYMIApUzWcAJn9ONjyQb2V
66w1Uehc1ZeFNkQAlGyoBydED83nd1ARdkYRv/22DCG0JzlNX9oM36Bs/mfm6KDp
YMCyOEZDEunG7CDmuSh4+Wd4OQJESS7H6EbouajXlZHWfjZUpcPfKrGfPZx719vR
fRMf9ci5a6Akfz956j5Tn6cetXQx6VF1jLciKnqDE8sd3Xx2CJxuHYj2MKivNSxq
hutEjGHhMaiswnIRQ0NNjGnq8QNfod3rHNHGa7rHL3UUdWSl8+TByh2XWH4fgTWk
rktdaDYJjXHW6TB8kP3+jZaSWat434f3AtEhmTfsFiGrBKiYawTrQyqtwSAe7cLY
2Yo1r6dTwUuiMB6ObZ/kS4wG7hL8jcmsgIwRYGHSzZ4aWEz6MmaAybJ6Dy66c6fR
D8DJxnPeOSzC1mIR2iKBpZ50ZUSosT3qtBLkhzP98EcWJtxyBVrt0Z9Xt8HwV0ae
0EuL27N7Hstmx7BeUmtM7z+mCNJ/iXUZsRbV2THHy+wS+p8ArvXYRClqAYjoexHl
1MOEJ0SoyBfPfIFPUn4EFW4K1qSqySO6Z7p13vtI2nFnNZ2J3wRcDwAI3fRlkorb
HeE2Vaieo7zFnh6zZQuMqriyJCPDeKlu62rlOj990lOM0UOdWzIUzCVO1/2dh+7l
JaXpKdxvLcWHqtbGTp6vOv+YsGYUzKkk01uNp+Oa3iDAJsJf3iZN0mZ0xPtQNPMX
HwFu7fDCYW1IP15zHUVnx/QU9YYVPnmO2MI9lQq8hrkiepO71LnFe194XEN4agVe
YNPW+svqMwvvlF6lGCrvkkT64YRKd+rMUeN7sbznLKL0uviTrmecKCLx7w1h5ro/
QmF58bagWysSzCU3jN9Ak6eoNyyCSVcfCyIBUdys8FRNaql1kZm+iQUSEis+3tTs
r/KBnnL60HgloS6UjRQyrmEr/eicaXua1Vf3ST/kp3v8CwYi6csz7Mx2OX6K4FhM
LmYwSN/XIAByGpS8OnoftQayL24+VdfIzrA8uXA/FH7YlqedduB22nXPyTBTI/Jw
sXcm7cdPCnXiV7mBc9tGs3CQA41H8aNrVKUababfFmyURniXicA50oxgNO5pEzyf
QfeC3pVmQs7JL5ESrUDOnq7mcuEtY2efTDEVPo3INYtF8ntft8VsIXMgjYvWtYow
ToA5nAtDgRr0p4gczBFbeKC3ATDfgfqmcd/vuX0SM5tRXGcfn8MX/Cv96KT/pvWy
XPt+18XF8aM9OkNZlaMUdSp00Mbu0QHxPEBYTwMtIKBg0jlV/OYg/gKEXlf9PlRL
lQNJCv65P9gLHU7MR44223sN2haguPIHxlZP5g/4uq4nw0z3T6L0Gwl12NeY7739
sE3GAVTMtzhfAi0eb68uNcbdTDkiTZMq9qeoGdXnW/R4+Ogh3mncF9Duh4HUasx/
7UnGJvx87Tc45pU4kvsPSgjRH60XJQwffJKw87Mg/Uj/WK/0CiZq85TQeKO5ixpx
alzJiGGJ5S95lLd8Ww/gq/gVZBlSHCB9IShDpcxgOe9W0dxoCmwMAeqYcWg0aFep
IXjwoKaGFiSNuP0pGCR5GocBBHq0Pm4gA6lTDluPoNuo6fdgllH+bV0+nLvp++WD
br3WDDvYnwJU0+IbtsTup5l4WZVaAsVxLdE8exCljFN21S3FIDGTdTpO/oIJ5umP
8xWoOyZ241oxGpp2pTfvXwUzG3hdHF+w2nIkrMGu18l87slBx6pn4UBP6lREuYG3
4zigQP/faW6HzVvkSyDEmyuMMrSg4sNzItgrZCQUVKINrxFFET0MuI0IHvFR9tv7
NRjjXPb8HsDQQXa5x7ahXx2gBCi98b+6phs7sNyGL2LE0l7lgOgU+u2aEuE6yVj6
v+uCmFCOnNC788syKanRSHduHr8CKhmj+cGoHWRz87j50J5INbSaQBvSZDF1ui2T
W6xzy4ZV1hJGhsveZ17uYlPq10Nt+VwMflcvymngtUau51lQpNMkWYji9mIdTYtM
AMuvYv9ANeW1wdExK7Rj73D8Coe9AdQElZ8O7SSPfTRcda/4sqBAsYElCM0dWFYw
RzgVIZ0udN6kbj0IezIovc7VB5PKWmUgcc5sujggh7awpAchJLMt9BZ3PQRCz2Pf
kaIrecemu8XHS79dKi1tv4F8qcS8xemMPY0DIH5xoyJWyjO9kuWDOTtMMplsk6f4
vinsXxk0rkiaDbmBXE6K8EvoZpNOfF07h615EbcZr0uUufefPHeqSaFB/8CpUGWg
bYWuKpvbSjtN37XAYpJQhYWfhdhBUy6K82bliKBaIiIUTRPMILwNqPnurVnI1lYT
7Ku+hx2Ulslas5finGCzLU4EUsbUNp6YLkweztGmStNkmC145jvEVXcpJe4XFstA
s/vTMiZcxJow2Zpe4USoAkLwuoRpr54zx/H0itIYubgo399xIOj3OkOiAoEJbDYB
WFRDmjqtBJDWYOerDIF3UShmCutu3uEsl/nLoAPkbjxjxYbyShgG5JQ/8BTg/nng
JQXqJjs1LHafzRxECWw9bDo2P6MU7Bn1RL64gLc8hxeCZnzvfJRd84iHUs0lmNkI
iBet9SrK6RDSX19DRqtiG5/3d+lBstGc7+8PmL2O7lHcr+0ffUIFrDR0IzRNmDV2
bvnnmvnHV3t2MI6UK2893c67WqX2JoGDzQ1ee/krhKgSQdyM8ZYIq0lYOaJ5xrMm
TSKuKQFZVwdRxTfw+K0S4xHLW8BGGhACUX9lnAumKH3w1HKUWqYinvYbrdJWMdk3
Kc4bGed7IuhLYTcBDHiyMEQapN3PYCIbmePw5Q9S9vTYOuiU73LoQg4xGVDXmzK0
b08dBDXX7Pw7n7l673z1n5bgqBRAvBDvkDI4z5sRoW3jMZpPTaMW4JT/KkbfzCGQ
77DPJqtP1OfQHM7iP5EmtfBmDswb1yxBmV5Cg71t6NSopsSzGDDOOcJuqR6Ty/ul
mkEcxszSJW/8AVeQMgUZQXPr6AOqsAkZKBg0btPoUZ6/EKxavCU/Zh9UscxJv7es
XmbdV+Oy7BZYnOIh7UXcxYtH5NiNzc2m3Hn3dCg730snX7joWIJlOK7qS2fKgHOe
fzk8bNH3QHXuXgQ5EMYU7EJzlhi7p01Arld54WZhiEzoBNOOSiN9ulc6u5PjwL5r
OoCMnYP4MSriRPx3f53epmwX/aawEe6Mn935OaZSJr+zCn4ZRcM+twjZsA69tqVg
EMaqZDfZ8ZVBVzCeoqzInsI93mebqC5BlTOv9OqKzxgHsE+JBfxcMydZOMGaIWiS
gqXg22bmm3t2EikuVkeOJWmFEZMpZizdBJ74LVTE9DxSqviJGL3Njvzobt4/U2wk
o5kSoFjiPKSh7jcAU9C+L1szUgcrQMlhrIJ7ccFktDQaHRaVLFzCJH3Vm6DbcFbL
5wXNOY7GkGKrklMP6WOTb0IJsLshDrH6twpvR1/aKFQTQVDtfdNrVukRVYO1IgM0
8l1I1+YdpOzkrgLwXGOPyIZuSzIxPmRpisPSk+Cr+72j0yaKPqapiXLECw43sp7u
h+obfiFFY9VBX2JMlFbsnB+BPIalUvIkFYmTBYEjD4woaTii7iJrKKQL2sDZarrL
1yyNcK5hV4nrEfOYvv5zUAAdXP77Wet0hlQ2YefumwrTFHPQRBvBhgKxRPgrypL/
tXE+eqON6jZA7Hr6QulycBKBIlAZtVYl3VqdeaFCQvlOY8C827pLgV6NkVn5iWER
vSFPYhvynlwpzrclYjkmdzR5x/EWVX3jyFmnU7K/gNAmn4tPBr+D3G77kRzd13dV
L8pal1JQfLiodf/x5tLM9pi9ISvaQFKpan6/ZlpzSvYQPLUaBnXHf/5oe7jpaHBL
7U7RBSN41hAgXdwgQNWPrOscyV8JTP9Cezzco/xEejvsmW3+wvAzqpPWY+c3XZAi
xWI7fsOEvosQ+kPA4EIfi16WUmcP2J1LkPtx+gUJh3ym7zm/m/CQmGxDdbNzpvg6
nddmidJTdqmfCc/SK0Gtg6OeOx8Z770RP0LDO7zWvja30Z1kEbopHOY0P28Dq17E
4tmaV/P58iHbPFiYIoZvKahByu/n8UG+8poQnF5yhTBs9YwpRiCOjX0ijlHn7KPN
6uRvLi7GeiVgP+lmai64aHwAbWdnyiLri4ERcxCPN7Gg19yzzWFFzD2uM+fiX/3b
u6H0uS/Ji0PZ3YHE35sHjgOeF9+ErF1E5ZW4rBTuAudHj8gAqExWPT3GIpx+BeFn
cB85Mnt9Zkcebeo2QRLw3i45t8xEpWV9UUGmtpZLkUJHUmB+Z+evXd0LdA5cvXNm
/U/VJyqAqSN8Urc0g1daTaAMFDxRjNxmJkI5RhXTzIBY29aTA3gjZfakOHeSzFJd
T06DEhoi5e+HPXBVTbP9ZqebNw1Hdm3sa+NTMIgWKfFRa+4nvS2GyFCYlboYxLRd
mQ4a4NHuaEdznzaBSBVeMxKZ0TH/7QJx7tI5EYbFpiVN1U3eMxhdEbA7jKWw/HZ5
sF6u8ggrmIo6sPYpLgmAhCklczrnruyJ+OxSCUc9+UJz97PCjGJmYpwvwmymlRn7
NFeLwyd5wsgjsd6fgcf/JCVSVOpMTbvOIVHkdGT47+l9v6Y18M3v8V/gAIldwaOA
/GA8x3nCsvHbNmbCJsgiBNjbijMPzi597quTyiI0/AMIdtCLJrcSI9F37YtCOOQ8
GZdO2zx6iWd8IsyqUNkqtsXowfagAgFsAbN7QeYPKRdfXbILy9B3C4CHjAlMEREW
8EyEPPXLm2+iuprvqcVXY/fnhC7kNNrZAsDfo/KYztPFGhjbJilwkCeoXh3nfwqi
NaWuP6dag9c3R+6o7l38SFdSKLT/qtu95qh3rk0gruEtnCdEWu8NYah1CgMS/xKZ
7M6JmUEwfSqO09dYDegqQG/366YBXCXXMwLXuF1caj+snGFULkcme98dfCz3Il9b
ZkgciEJ6enrUm7K/w+dEpFXDnpZHwfBEJUJGUd433tbWVun8+kY25krzoAxFGv8C
mJR8GbVBxVb4PRkkTPMcUf5VgOm65R6/aC/y8Vz2ifheB6KdckWF0PhhUAJvUSqK
JDwOEiF8O3HRwVJYXrYP/gDg1bdRXyNund+3/ADH57wKHORKYndX2v+zUmfb5cLY
NZ6kFbdm1PBV7bL2n6DhlrSkHia2LBfxWCt4Q+HuvPeyXKLE+zcBSqt6q8dIsRCl
oDGHmrMHBBtG+zffnRZNeFXZ6mj9wjssTcdd7uM3JskJBbAGzRtDt8loTykC33Pd
M7vw2dLxr7ZmStSaGn5W48hG3Gc+0A3buILbZM6g3IJf1rKoLATym81J8sfv1K/T
vCxUGFUl1avRdHIEhlpA0VNem35BpCAQ6KMEx0Bdc6awvSfbGnZwKshQSAHrmOZY
Dunn7E0QjFbT9E7/4er52MEeKR3avlZVRua4A/4VxgWwMtkdVAVwdPYn2P7djKvz
WGU96qY19vlI8zS+1jZkBv9iUEN3DRSmm6I9uG6i/gkV3H5AoQaDt6B16KlWgBJb
KnL86NLmvjtUqBxuCNQ+KATRFLhCKbVbyb0+XFT38U008UBlll1cCJp370MbYNPc
nzLtvkBxwcaEClQV/kDt9Z3tZvRKT8AyQl6V9o4KKnrYjxdOO0gDtTaoeTLDlWF8
N6GxKLAaC97AIOdi1CWAq+G0krcEf6ulHiIihfV6GsV/M1hVM5j0G/sJ8L4aJr40
eIyFtiILfiVuIzKNPIMR94tTxqF13I2RueMQdWXkOFthLBMC7peDT7PyN2j5QAiu
em9OW0kT1LdnKHcSRrO/8Uqr5uoU6Rcu+7Qm+ImFRe9PB0SSSMUAvY1mUDt4qmOX
qAzH+scQVpNfwEtOfymH0mQ+lZfHc8aKog860FywCa1zNO1BI1CGHyWJSfGvcCgn
Z8sNzfPUri+98J10wZqfyaBzsCNXjk9O1C11xuB6QRvn1CgqLak2MMiPIAlv5Ufc
qnMyQFvOSvqJ6+aEhTDbk67/ig8V1ggrb1d1icc+qCqdX9+faIZMqqSUbOh11LPK
/SemoeSesoMmVmXCIIxjfwZeG+qL3r3GCoZlsL/q0EcguOS+Oe3AnG/gcBbGJ1Hs
qdOCAWtKBs2gimtTQ6Iigwy1W8eidTEewFj/ZeducoBjnpYl/yOmZCwXuDDr27oy
mWDSBMuMi8JL1siBQZsIyYbIP21pHM1DIFPl4OkrYB4JSpk4tm5WWClRr0NZm3uE
mYpmSBYfxnTuI7bMjPCK7V+K1Wj+nit4VsA+tsiiPRQEgzpG3wbqjWGaaitcb4a4
tpnpk1kfAsIjvUWto7Z4npQytzJPZCInYPMq6JYjcr8K/cT+KHMrKRYaZknkOcoc
MieSnhBHATLx4+leyI09dtXUIJyQQNq1h0OAnskGSSXSLxQ+ru3w829ANQ55QL0g
TalgG91xdJ5nwwjDYnp07kOWWbjUS8zCLJUGvDutHr5unG/XOFAMDXQOiF4CATjb
W6D/xCbpN+dhhXmApYVFbY8GS6XOlEFxCOoN6MSw7RDCHOIykgXWVIEhNHAKRiD6
l6/RPpx1UvWmfJXcavGDdK+mlEye4aXiOTdE7gBti7AfCOEKVsAGsUO84W+XEbeM
ZQvjX0vWS/jIhGIjpghOvAV1TDr3PEdcZ1fmHyX3SG71paW7+ddW5fIoCgDeOLi6
a5l+4iGQkAhZcFYB91Bl2WA1pmVNQWhXgHKYssqpcfudZI7i64y34dNgYQNXmNlm
UKSJT//tTmdLodZJfATjUWfr06xKICaLHtjJ7u2BdQezK3ePFPgvfaLYZKyxnmTD
F4GBBrq06GYAPVw/f4ghzxsLJZMo5xygvi562fGlvGiie5edIoJsH1Q8PlgLJcGF
/2Li2hbFH3ca2cCpw0f9iyBSPtlOmyW0jY7j//tRzoZfVdttEWaiZEQjeAxdc04L
Wm4K83WO9MzRaXa3IptOLceZHlTssuT9uyun60ZrzQQ+Eok95ah+XGwk9m6ygR/O
YFCqISZm0STBNHPLjaL+BZ3mn0bkkpKjnEyHQT+LgLiiOk9o1fSvVf2hOwfAUCBu
9TpGlCVrJIiX0+0aAMd2P5GJsKlVU0Z6QR16RUZZDeaaomPRVQOGiKMvf5EgdFSj
Sv9iTarpG2vTgs7peu1HeBXjWuLuWYXg1/D0WghIi8FfTIK6BYlZZYDF8nfBa7D+
QI2Hg4eftSbDjmE0O//BrFEC4IRUflu7xzAWreU5eHsBTyTXzMirMy+EBFyLCiAn
12e7sB36wHYDjo12KuUSfOMUJ/RRbQ1xlxM+OsyrGel3qCpLBcnufWys6EQnJsvL
mLwA0fe45zz+cX4Yqm7jHwg0rWnD23clIDicpSWeSrZSiqLaMlHEq0qVH0G1Vg4x
hBS9ww0fMv7jaQkl4b/P3TAmdP61hweehMEZoxxoOfa60qEis1jdblJpqXWki/p2
PYhCLwyLUKDscV9Wk9ETCyce4d4qYDJsiqwNJ/kCNih4WrOZJXsiPucx222DN7SO
5WvjA38DVsCUAnJKM4RzH1CKRp8Z6xJ/cOyj2QZJND2oZ5sG/lGEHVa39pvNhP95
KmHDasGmy5pWIE2eerfJBeo+nH33/QCNCFBTQ+E52NliDnsjoZrJ/0PrdmCi+NXx
wefD7zaML2u1/y2u3AAlSrrvrY0VuKIH1nCpSYqrTzrS5ihzIpsogtK6YyXjbdzM
KOjfoSBMR/48Vflbxq18qxnS1Da/32DaG5wamAhSodoGJmlHZRrChp2rcBuf30SI
90K2a0hJyHfh547Dl9wjC1opiu+dzZah5IMqpTS9LU+Ts3H5nm3I9EuqpBJea/F3
1F4YoeUNl+/mCzH7SLmFk5OyJPnc00m7a7DKC2lyJ9zFnfzOp4alM9IRY1qDmMhS
M6acmbaCHf2v+cGelVeJuNqJOpbMSDec0cvvQQUZAkXHJTiyAkfrc19fe6pu4EsV
X76CUH/LaymVpV11ipeB3dgYCHOSMLWxYm9c7GA2V/k1vDopQspPITkuKKrl2Q3n
cDjG3ue5+wwqXYlP7V/YtlkHw32rpi3wQR5nU4kAwtGqmvh5tJrSHjK7HKeXNlnr
zyXJaCoIzzAVaEZeFZMYDWlA3MzOZ+TlWelmq/mdjmxejvugTva8Vnjuc581Locf
VQiFILBswraCJW2Bxo1g3y608pCR+vQGwPwotMZv1T1lfhv2wGfOmnym8rOdZYYz
OdR3FkrWHdwU98XEnFoGSkGtBDXwPVwWnS0lIv7tMIomxP6H49IJiwKUK4K0ra6o
apk5fDqfU4nVriBgyqozF+5d/3iI2LC1dpeqRvXawZXtR7wNdaI5cMmoRThK4mvk
Kemhfg+K+EcFvFQp79OGDQV3zH74BEp3/RNg84XYU5i915Z393jzQ3vjTFCtXqvg
L+0krwLt6JdxtrQwz0mqFtbSvnQAHBN0s3g/wCYXC6uqHp1gAxOo9UMkeP2jjPBk
Minru1+FOZ3xR2v7NRMWBlP45MtAs2a5+MGMGj4dPdYKDUFvfi1FV++l/eGsxDGL
wrSA484Fr14YTNPnRxKrRd2iZryvbKD9Iq3ZrvXq4k5N4Ludn87x9WkCuzF0OISR
9sHssKVAalLRbhNDtgPJ8BJm3eWhxdV4iO1QBAcaUOXDiGNGD8lmsMWTxMmdsC4I
bDDrTlrYGWkEfZ/K6LbQiBvss6oquV/+W+AHOUsw2KXInaLVEHE36xKxkkKZWgM0
TfLpjYxn1dtB1nyc8huO3w6czPACux+HXN5+azpvGJXxMaRI66jdjLwqbirWEZ0v
QDM0HsX5Stgz+H/wAcCLtT8wI8ZhggLiu6w6Zgm8lhAO1epSFt88D8nJstChITGg
+QQuzH3I3YMvDHKsdyKIa+3eU7b5kCAgilYB09612FNShs7mss5q3jLimT9IJiXI
miRumMAhYXriQ08bQmZOOEWHmpjdTbBjPTovTdpXCHEnc23ZY7xQXqc2by66AgLD
AR/cEg2gAnP61mkXo8+01QeCQc0T7Egwc3/a5Q1f6P35fVTbwTdC0QbE5XMuwenO
iWBZF0jmKqSHbtF1GJ6gQVqfWU+U3KU/Pfc62G3OQ/NGZIKQFWAYTOq2scqDrcNb
IlOtBg/GuPeDriayuaHPoV+z7/q9OZfmiRR7kKgKZZ7ASyk1BEOAXh8zha2A4kDy
nlL4eZYPvLo3K06gxC7J/NTMZbN3nQQ90JS06IGp0u8/Zt5Gv/kNEsmoDa9ypEhr
8kY63HVto1wivgN9xw4b7e5SA2rAaDYTaLBdrIfpNT9gWYT97PsmdAfLiK7Vp0d5
nxo0enBJvdZvmuA/1oU68RO1UDkdO7zvlJ03+smpDgDgBaWRzyctG9Gvgc1nAZlU
F4mGTu6FY+3AG5quyWhsnJb5AZwtiwtUpgNU++oZPx877GC7HHL4EcwIpgwlZjkY
ag2P0ZgffiELbbdPN4LbFJWwtIIRJVhwa6YR9yVWTwgWNOvWbbmEYFyT3nM50I5R
OlA0P8A9x5WwzfgzGBZbRTT60+J8vHh9PcsJwZX7iuArkJHxLhcf+CCP4sIiKaNH
IIVWVwym8HEfF/tWcRwTXF26yWZ0HPdpopfICQAB06wdAsHChcKTPcsFW3YcAyif
vpKc9gGVI92RtTQZ8I9zZ603TsWylzJfyAQ8AiPuyeV8wYatuPA7E97n4BZSgc8a
FBAyyHz4a6izI6HstVLhl9QFjzuHjPrAqenKjFdoxNYFl2m7iS57E7hxjDDodqT8
MCVl+bV0lUn9mtwW7X12uD/VTYx3vhcGOUaL2+iCYRT9rIONpugKwyVOwd+mTRui
CUKWFVa5chbShg4S7rKNpEPrNOY8LBdzJSjGmEARXku+1mZXB+h1a63UkLYZmFhM
wtlJWIerafiZa/AT1h62MCuoOJxtE9aNvQnXUUtVCPpt83K0Tip++Mb1gIIQQzpH
HoJLxBUo4VNvvLFBmDvZUhZpPpatzjTfiuzwhEMil0ValhlKGJWSITJn09hvpEhb
X5no7fPMg7MDkRi1D5h+k1IjY1QvJTMD8PbRH8R2WYbjMAxfwGwOI94uz7tNsqC/
EzjR1+EkdaIKxqnMkoEXoGJqaYXDQIbbhJteq7J5VYSmIwwKv0zQSMrRwHE9dRzP
ypkzgYM/1sHTyJECu91LNwOnhOHXekvvrVdA14s4To3cy5cm3PUGCbBDb7WIX5Gq
T7u/xXqczHfsFxOvksrnvO3NjCjHXBBP+9K6gRLJ4qz32Cpx7b1p0TN+8Co2UHW/
kQSFEcw73quEjUdBQOL02nw6JGeZj1mmHlQU8XmZ8GTjzFdcLKSO+ZXY49I/UeRz
828hLqYE01izR0uMR8xE/wRSM0yRgz6WgqfyWoLP2JgL++6f0UJeEddDng0oxSog
sKqZ3Y5xI1VDJn1nwv1J0E2r9axsCtc/7Pm9EZsID+je6tbZup5ANw8mGNtDqQYL
6YDOvN3rpoLI56Ke1jrKevaK9N9x6eV7QW3dRdGX9MIdU/X4ZZH9CruA0RlW9r0n
pNcRv5Whhy2JzTjszsN4bKgOWZ6k4feG3YIQpPFwJU/Ux4uqcDZn+VU2F0E0xvsE
OutWdfs/NU2apOqhDOaJFpqH32G6vTvbf9fl0rDMCAa7dIA5I5UFXDGR5HAaKC1u
o2ce7POs1U4Dyj0T/qIY2/Bbr+6twplMSXp9K0qm2BYvmwvMZF46bHWxxfg9LG/B
1q2nn4zNUecNbY17R+52VgR51lgYYauiPaoi8SCI3c/py4fdn3vb2nlONsuZ7oEt
z35zQ8K+ZRNYkwIkbZ21mlPAin8NEjo1fqK3ZoVeleZ+eHStYHCaWxsUiXgjuPQD
3LyBo3SMU9jP+oDrQctN3kmLe0e3LE7tVx056VqKg8H3ChLPrs3OhWoXa+x9H8Nj
JIyAnZQxD+U3GREuAtweteJUtYXT0Bf0fG/iW6KC3Ya3UtqvkE9eqshtwVUjEzCy
4Si9qlurwCcK5x1zE0iGzkLILLuM/H0QpZGxiIHN3qkUtPWKqGPlRNU7TRS7P0H2
Y7Jg6ydqOZ/q62zCUQ+eFdhCDYpwTtPXftyKSqRQ7JPkVIeR6XPrqy55dd7p2BOl
Vvqt0k0KIJD9W1w+fdlju+bMXquInw8c7qC9dhoICAurmbcm/Q5MXffGvDoEq9qQ
N5Yw/JQF8D4UAnPHg06egnyKzoD9950VEEU/HNHmncLE8TFPw5WCNOeD6QIVjnh/
Wb9Js77qAKwNPZBhpiqw6ZESWJhMJgUWoN4SYa3gCKLAnsE7IEuUS8VMmVwxSSg2
eeIAX1erSlOQN1KH1GvzLKdLwVNrWkugu5u6RbWwFGPuKfNQAme30sk1AfSyXFL2
d99TW0+OsX0fP54QWr5Ijr2FhbLWgbQ5irJHcjA5J6bV6eQfD0LzFZl2Zs8RYBae
uQpsE3VTgQ56eJgqHBAkNgDd5SzkF5DCOeymfqitmEYgpSW+nZo12OqaaQideBLu
IGmxAE71RbGkMFtDDjA+6O27zD5m3R9Lgaz7eev4lqFYEZhNjM83vG7OlXk/xSb5
8a2PkYPO/YHZsu6D0IHC21QCpUIevEQKyttWxHvpo629qDMl1uf7h4lLysbFO21+
IFJwEZ9WlO+3VYB0QP9dBklcnE6WC9HmHtztxbs7c6Nh5WkddT+Qc1uhjC6jySlp
Q6mUgg4uQsQA2fbKFLC5lSrh97GXb7WR5PhIhMXuMHdTYlHo1hWlIBcr7TSDAGoD
iKsCt84Y8ub1M+opvMXS+0s9YukI+QmmJu1LitqfaVYMXI37ud8M3K1FTk4pI/J5
/c/MVcntBVYFUmTzWJKO+zxmMIt5ehIKe31PoylOcqZd9A15WnYAmntqXWZG4FBK
xEUEpOB8sewZuINYAkqyqiIxHXZT258/bCt7OLiDduvgNVY3WIi7CUkXQjzVkSrT
nbUCuMoeiScfCC/2wty+3ma70u7FsNKLLoH3ikHW/YNUB8//J45qSRR24y4uhWuJ
vcHpRkQ+mdPLniRUpsAlux+xXlU55a58Wqe8KbKRi4svBqEYMQYybITH0t8S9eOl
d1ECyV+nxdZxGz8HlI3xjy2WIIM/PtRMsVmFe6Kn/iHDycQoTRpiIn+X3mrJwlks
PbFnSCJk/eB/e3cWCpyrUIF2grskdSGteS9P6/Kv7tdRJEMvxj8NEcX3/nfwdTo6
zvQz1YvkbZk6qpXSQfNyC/SgZwJuU4S1Aotm4kfJ2kkYQXWTCq96li6JqpOdTJOv
cuwVFjy4cTh7/Wzgv2SpvQzZbrUa/6BGh/VQtpcsZk+hTYD/IObW1YV7dWLkjIv1
Wo+PngvRiyzdMoXWWcFBHLnI65C5U9WVySuEZTppvwt6i15dU3ncob8rGibFzhCN
Ck6+GSY+0p0qanid2LM7yl7MXXSkTcAQDuM/bae4X/r7X2466r3qMeEwchbd2Mf/
aHX5dCk++HVqm3oqoqZ2RzAVO2lUmcE59U+QuB1b2wYK3mR1e9ovlGx0QTilq02E
gcst106DmdcIyZ/kU057S0ZHT1eExrjdDNGWnnEO3ktvM+ECZWrEX6DBZDLINVZq
iB+zD5jAjEscAn4hFvnUWSiEKAUkjBkuV98F25r5mlislcAstA21Wgth4WCoumSN
UI035tUJuE882aYrvi1MNNP6nXV95orj+b5uLkyVHLUAZNZbPF+K0zRR7xT7Xz72
3CUhDO7kL+riLbc+c3Xt0dDCLtG5WuOFpB4l6c/sq2ggT/l1+h0UgFTG9c4nOKCT
1Pw/qqehpeS/8KbDCFb4+TTSgk5nzWHJ1xAg6W1+GiiKPUXERWN9IgEJLmhC0sEH
xsFVTuEJUnM0uDseYCobLDKmkczbTBW/aqCh96+IHAmxDQnX0VPQiDL+BRIkowDa
8p+puKDQNWV2CfCoOSzyYiP0IOTVe4RCP9ejPR3ImwSv8yEKrwBIKAjwqRN2eEgS
KEc/F9MtdbsNqSV3VjiOVotI3T8IY4kxJUo3Q08CRdf6Y+PoM3iZ66gYWdWxR6YU
O7ExQrHzyvif7pTawLsJkqF29mcVaG+NjmaU6Xh4tPT2qj+tsuSojw8mjTHbgRAZ
azXhNVmPsybOToSDj6Rk93lrinxjYdtimvQQRCmeeEyo1dXJgzCACUhwXIHZrlCF
oKJ/9X4gyQ8x0yhAca1W9tcWu99qJuOGlV3TQWIqXn8kemRKfwbXAAr2KUrO9C6x
BqBBMMHOfE8YDOOYfWR1/ptmd1b8W+xXCb5EyOBZV/nV01VF7lcUzQn0h3Nz3iYj
//Es2BRx0RQ80tdKylO/gClqwXn8A8nZzt+PllyR8/UfNur9rioNZbvxRYnvbQEJ
tTp/XSoh1USFpqJNP5VHVrW8fiWcoIugI5StM/5uCDxd/4Jd0sAbwFpKKLJ+EXJa
QSpjHfaH01Z9Ve5/HCOLBWKl1bd4cnlP5a+9Lr/iWuZQpkVYmRqGaRBVdJm2FJay
1oZvbbbR5OVvE/wmSy+Otr2tHPpf2/RgWPk1wdSmjMOsVsVyaoXf2IgR8HTFuTZL
65te5WZXgAxaNTjvuwQN/b26RR++FDlghChKK+niaCzWhFr3qHIbYa06+8zlqX97
l+MSkjJIgCFMKdfzxAlh7q/C5zVRy4eOYVrBOLNYq7Ito+B5KWXQU0/iITv90ZnA
kg7+b4HZMYt1emprCmYC5zwzvbdFencUbDulwdCA/uFTRDxzzoRazPU8dUrU424B
IdFf6GJ6UfaiijFdj1GguDKEUbubhczz0Wuj59av/lc94lh7AltR1BgaO0ptJ4z8
v4jwICNZ5wGM6PALOAT7KntwfPR00+Jhx4ciUuUkzdC8MMoCPYLz4xIDeKWedKFM
+mtLn87ADYuB2SpsFfq2L7dYuab/NZj8wEPmOiS7AnjpHmU3h8fOm8pcXiKS6Z6d
0OTYte6qNF9Rm/XXy7jo9OM2MZJ8m4xYn44c+8Sl/2nBwtur14y605LPLfO75usk
LUprU92nSkZ334f09PLy1ytm2GSTallBXflKl37m1ITS3ualYyjqGdRT5uS/anj2
G51onenRzCy8uUIiwqjXC6+R4pOY7kP/luRgcjRW6M3/xh/DvnNX3I5ayjZ7lJU/
+IGM9FGLEHsg0lvVCAeKhzWHx4Cq2Hc82n0vz3XDWDRofxV2lotx/ZTtcaOJe72f
WODRy9e9yqKerRb7B7lYsk6oSMZSEe8WBgOwTbD88OlZ0buQeY6dxp5hprcelEeW
iuidHiV41rCid8XaevM1znWBCckSDA2GeRBZHQR7NX65/uvobwH0FNlesM7tBalC
uANOQFlp20RyXVIQK12+t2ecRJR4UbazyHdDlt3eQPjbmcK0pxK2Au5bJF8Pnm0V
YhP1vRs1BbE6YssomDpja74U6nTgUKOjBFxn8AgJdDVLRpFhtbqfScdT0UxXyhFA
y+My7FBx+Rv/xbzWZLFXOTN+chYUMjf6jytt+Qq8+kbYk38oRfLvojySm1BWXD9P
UBnUHey/x9D5Ju0kx8LOlyb1DkHgblUz8VFIrLBOT9b5T4UHpSOj7x6iqo1T4EXv
pVL+TY7VRdRk988A9X6tlq1IKR/sCuibzty8zT4a3i3ITFZp/fwYQTDtB/IsNW9W
L3gG7vyHws6Brnmcmpsv4LB92cnsUOpewIz8H3qxSR+J748IDV8+cOVnfLRrxfrB
BETCPp9Kj8467iD+xFtddxPBm50xYPr8t7Ul/Ybt8I24lSyr+nc/q+fTth9vzUHe
xHO1Ok2USSIdduNHBn3K4nWMc97l0+Dx0GEz7G+xz7zjYIrKBWm5IU4m/4Mtgt7/
V+BtcmTuBvYpYL7z8xbGOb2+jMKgb6TaOXun1aE5LI78KrN4PoADh/Zb+rtbPGGu
nKYdL3KPNAjg5xSfpouvtqR/nOEo5rv7uXmyHyoXH69GeZwV6ySDwxznBZhHKFpp
//OJRUQpOYC0DKqWwpJAxv5kXeCrosqxG5Tmk6kA+hHkd83aNrwtzTHbYUmn1X9Q
fWorBFmdbvMg56zqdhZDEom0WvtuC/zOlRGLv6EMqbLU42+fe5JLSVLBbUbu3oYE
bKIaj4kp9Yqr/gQFpRj0xh0A/I8n+MHz2JQuodwDOgAchUo317ZZ1n1U690rPAlq
DcqvJLkvYrF22v9MMeF6LfyxQB8wwMO+WaF/QA3I0M14g4Zu1KQMh6vpPGAgZWLi
EKokRjZAOTmPKEOzJ0D/N81TsCqSLP3qY4LBTNMLDdCmPPmhXq1lFtGAsVVIcbzc
4d2cIvkTx/CQycXe3gyFte9G8E0P3OFIGBGQyW18cAuDWuZUnR6iNhlFDZwbFGnf
3Fub9shryDe1jL3BFp8OCzQQje+rM9efl8NF+Y0Rwsk40zEH5FlWSYqHhyYvZG1o
BGzg6DeeH9gsipP5r3fA4n/TirjH2Vc5UgXFM9rv49ptBKjenUTnOhxhO9d2ZkAy
0aKN4gJlm1wY4pyAPhzHf/0ExRgs44FwrpBRVrNysuXaoWCKEJPQTjUUiN/1vT9I
qzahzOcEwN3i6PQKQ4DJoCLckOiDY0Tffom7DujUfdqzbxi13DOZB1HFJiFHH+EJ
OlSjmM/bF7/XURNcQaWn9pQ3bXRvV908pF+O3TbEe6al4O2PlXqHg2oAw2jixJEX
ID2xqVslaCKoeH8A8YqyIo2l5Dp5ka5+1f4ZJnX6MnD5nwnxksMEeqVGBdr3rVSK
TenB4JlvpuA7/3euzm24irCBrXNxnKkOW2nVEzfB8xk3JVAEd4gg4npVQPK86LBT
uHaT1PK4ooeEJrXma91jNOXkmsHqyWYZuOiY9uhH0j+bjJFzKrDHDEpCQfW+zU2H
EYqIjakvHUwZsliv9/6oxw+LjZp1knSCXXVWP/RPGMdA9q9GEmhnncc8zJbrkMzJ
kpwJ5brf7mCFxB0Ctiv8wVByJqUIMntNnNt3I1F+qQ8qHT7/97gDjxmim8Rp1YP5
LVuuz63y8L9OxVWN3Dm5AyOaUpK3jeSjVgrfx9JwNidclF504AxdLKGdnZxjal+8
1scZEZutqQRbBH3vEOr+/1CFSsTRO4SvMEFv0jqR0va7erVkM4LwEJULvi4VLRW1
wrX+O3CRN4o++walvMTfFK3dRyuGurzAYS3yBoW7dUA5QOSQIpTLPK1wjNmpAWFa
HFZ4zn4g3JN2HEDZ8qg+b4uNiIXno4N3Wgt9h1EL6ycyn1vBoG6egmGZ16urWms7
Oc6mJkjDJ17vrYnQYe090ZrdWYVmpX0Qym9drKR0tRXxqKBlcVqm0QmzNdcDWIdK
1uYWKGvAS27iR4QAkC0TA35U/PqTfBqyMnxNk+POjbWulXQZYIgXsUseMkasba9V
zBLBG+gnvlLFaHrX51xiW51M3k8UeABBU7DJrR8kh6uX4rzKkDcuYoF+JtUP66GX
llkrXWjwJxldl6chPc5Q6rn0uKsTeOV79aMT6/d67Tg+QvAm8fh9gi7GlnPogzs5
1kU6COEbNPn8QsAZkVDb7gY2hZFhGC7UgPIpFa+gJfiPzpyE4bNXDp0tCjTESPCy
MTVYBX3Lmrv42PXjDD8Gu/nSm8Yo9crCO5Hsu484myXPRgaQNWeZu6ThiTOYyQTl
TjnRy0Rjkzj22ZPrGXFy7naLmkX4cZzmA2V4ZidL9yruXoP+O3stzv4G9tNW3W8i
ErV0UjGlWBquGFbjs8KzTF7ipr7WTkEg3IEHGB+W0BfCF2wh8GRu15nS/By8extR
Xct1r1mzegCfGeUKM6paQ9V8hBTIAgyxsRW8K5gMc7SYXzadKx4THJQIo6RgPNXu
049Um+3KwXDRaqaAGoL0Uf10cTAT2lo8hea6Hs8BUEIe81DzdDLdkeATuU4c/1js
nGUJfsRDMwE5NsJES7NAmE6DWxE+VNkDBDP2NApzL1G/RwxFGv3I8/m/w/lejPv1
z6WXig6zcGjSdNzvTs9/RT/zwzp61AaQ6m4Zwj9QRfY2YxndI0vT5gjife/Sluwy
GGRsI6y71awRkE7/OCqjsLrYRqD6bqlc7mpRrm7G4BHTbKECTpBkFMO5hiYMJC2o
zOz9kGvEy1z9gboBP3SaJj3QlhsnO/LcRBAr8BsS4SUm0Epsj21wProLAaJq5E32
ugfmqOfK2ao6/DVtIzicJRzox9CRtTgTTlZ1GtkCo3mXon9cuCILXVIyIpmkBE4Q
A3dLpA1pXQaKpVDrWIYoOPiTAQM75KRCWN9RAgQkqn7/P7ZOlAcLiSRlJQo2Vovl
5BPC5iKvMmmwvWhTdLqnoYlWFgxJ45v5rnxfGyJ9vAZq03FlaRlQabVsQ90nflcC
yDRlWRqx6kGsUCLfpLZOwd8n6LAyJwcMvChgUuWqw4FQbisMr+pOQjoxblS1JvED
4/I8maey9ak0ifT0FoDZhbOEe4QZZ8ctBu54neiFnYy07TQUk08b3J0lWO9YlnDL
dkEp61aGaE8H21MdMxwdHgs3wjVO/Ca4M2YVLEicyWddb5L5KvZnx7WWFxVqWXox
lyVNmYaZc+1uA04eTQxUwRhy6CCFQtvxa5xQjXF95JmLWvepmXkgi8q05Bxyq3JZ
LZiTrfMtPndwGT4pMfm7rK4pSmdZfBFMxzIkkqRaaAh9rPntbM62Op9g+jBxRPnX
oqI5bjep9DNlUPWiiewbJvwU4LsAlsihgfCYcRCUPKFnYPu6/U2hczX1PnUmAiZl
/BVidPm5vXbw7NEbOaVN4KtMY+QFvWmok1OVgJLVz4mgO5ID/9AInOwoTE8E+n+R
yD5zqQRZtrKB3xN22SNCz11PxwCLMvcZhf2SZ410uVZBtcgiAdVco+RD4lt1y6pF
ZFdAylZxBmB3yQHZ8vqeg244ApH4Q15AYSYtMKaj/9EzBKFCR5Joi0Stlu7xKmzf
4Hh1fwtHExbMtmn4vzc+bfI0sbkWv8y8T34L5huP+Zl6hMZgzBLZgRZfV2h1Ette
KGPc1/LK12YNBZCoY4cxCX6Bqg30RfucLOiR0DYj8K/CW93pmN0IxVHBnwsXj1mj
P8IpIb6eFof6kYGAu6mDedcocFWklGOOVfeNUzOZrj0AQJL85trKl8w3QIXLqYPD
hyTsVTzcze7CfdBYVSuW5sg1PfFMqeBR5DFwxZKD7wXDbOeHTB/sLl+C4RVlMk1T
T1AtxSsurU841M5DNNIZHZjXn2kBNeDCo6OeD3ABZ+NHttDa+JofQl/zLQHWepl3
z8xUalvAjjvgz2apPMizlDo5NnnEPn8FhcKXK+7snMBPnUu73RHSxoa4sSuhn3VI
VStAbtB8piPmz5GT13qYTCiBxjGC0/1IwxIbPr/2/zYapV8N42HXm8Z39lSq00gO
unNAoeX1Eck1Xga4L+ZWtnBkYww49luA2dSmqnj7oDiIxCd7u3LebIcqt3N75fWm
w5Pupl8xomkQQymiqGSpA1aKzBPn9RqIqxHQfvvcKkn2c8NdPlbsphayGKNtIOHG
hLL+hDlBIkCUQ7oyE205gkgYHrpKWst+hexFYVEy2yVV9PXSVp2CmpHhX70oUGFK
IKy5SujmbV0xPs5lbhfaaooCMVxaOxzL/U2yXBF2cb5bQnLWhNUB0hAqRZvYLSo5
oMzRjwT1DvD+YQESy92elFQDs++PzNqgnC3AbjYLWdkzHUlc+yatfo0OJKBgjJyN
MY3LBDA+wj7S33xgKRQhJGoPvT6dsgLIkkkGfpQHFBZ6O7s4D3yYkkIW3rHhkoj5
2vBIbq4ixG4lQ+AJjagIGhqNTOUoLDY4fHsoFFUj46+utAWeop9ipFW4XwTWMRre
k8AAWMFEKwMKTZRQAb8NImF3O8JlA0TKQ7EzLGzrnwkjyIpJoo6hT6QD4NPoQ344
+t6yGbz/AnlLmHAaHhBdLZwHiyGVKUBZSarSe1jbBz3JYlXMu4zOPqhh0r1Pvnh/
l3bSHAC7rRs7eYW6pLi+msVMJsyI5lRWbe16QaLMe0cSX6GwAld6qOh6LAnb91e+
nUjsTtN4oxxH7RoTngJQncm6oRFkAXQySPLFLh4ZBR06O64qHuRqumwssVbuQjxG
wL7HrcMxEdv9H3EGQfKUmH4a0AwZcycvEeyJHsA2AerBhZvWG2e/J2AoSnx04gBd
E0wXeL6SAElJZKykv1o3+fxIone8PUOkZzhaNuNClvSG0FeF9XlG4YrFU8GRu+fE
RVXYuZCNcPFXUWupoHJCXYqxrry+FpAxKdiYJ3O0HdW9zpLcQlVDmNCqv9yXCHPt
Wh2nXMANVHa16Yu2glBQbdOfdcstBsCIK2bYlNWmqMiZ3vE0k2VRh2M+vUQjGV7U
03ZRh5CUPSobec//O3/0o7WQsYAvyMN3tKxhCMC00LqZBkfh9MNhclHy7Yv26Zm/
d/P1KcMWv0QYZa0Nl4p331S2lQYiY8OxhmybwX2jriymbajxdW2sSqCFNeWhiR83
dKKp3tDCb65Ae1tYIyVjK8QnH+R52qmsx3AdjUrfkS+XtpmMnfoH3OKtYyfMO/j9
A/3t7Z7/WlQlps29fUe2C8OTOBEHh25ZfnPlbAt4iekoauNMCGrwb8g8RJcwOzpE
+sYStwuuVlrLlz++0UzYhRPDX75Dth6OMRuGmtjbotsvUobs3KM1pfZdQZx2n1x9
Hb8dvzDZp0Hc8oxorn1MVT+nzh64k+ArY1odhs1ksRHLVp0vKVMMGuC0DAmY0y4U
y2RDT4I3rYocldxwKSW8I02Mq4f3MMTfydYEhqHHVC3GUe7hUfdMQ7vXIuKJsFKq
3M1ayzsfkDk+tDrTEzrep4UscX2rvE5mjhwUYFu8N2ZzQrVOeHk7sZxmAzB3ylED
YRPpN7mCvvC7PAx+AzL3fiRxHvsYJOFU5kAkJz20afegFAvPCS2XWjYYFUIr88ua
djP6i4E9SuZ7jFB/AoqufbX8+BBrHijsc87K3zScGwHfDjyTVutwavSNHcGFs4Tn
k3snHhExEzCneprlt8mSc65GyGzQftug9zos0kapM2XN9cv51rLZGrjrvo8z2Ht1
F74UZfRmrbegNv37qtk5Yfsl+yo7MbjPn9vr7HRVTBSEyz6rok5bE+/1AKJAT6at
3A5HemAVb6k7115yEoyAoKberDHXKr7AWeSaT3Xi9bt+K1uq+vIMeJZmculoXrz/
VxKi05OiKzjra+Mfqd+yt9Ww4CwlNiYVR9DtUqDN4tA9TmYdh3biQcw/+hvT9i1w
tPjrJwE18JuaC8ae7enjrXx4L2x13VTZSJhCJoxpH2KgsV3F7vE+Xfs3LG0k1t2Z
/gtaHU0g2yADNPp6rL+3/dcZjtBDmrnsrXdHa3KVAv7V74DbCLZSxAWsbMy7I/7c
IOTThNUjPPflsM7lqeBiiArIrbcGR2DTnbzn1j9z7RjJXObeDgI7xHPSbQherTEt
+64i462emcTEfoBRXJ+ZSIGHcIbpguVhcM5yHFyfWhvLNmefQq0oaBHNh7B79yn4
m3aa2WlGaHAonBK1fhgLEWEDWfiyGL1DojboOjiF/i2fMvpXwJ/n6eTWYTowByqH
nvOeWYtCP21ZbrWKiI/MoIHBAo94toUx3uqnMQPJY0B5ax/pxemoXsIPBNcbNmdd
32nzMo0MtmU/maXLZUHIIs0+g4N+Wj6mpJYv20gqAFI0+LeVkjQx33ZhvxkcsOCv
FUbE54/veAVbNg8sc7yq+AKT4+hVOeV+JwTdZNHEBA9JiL6UA3noyobjXyP3kq2/
APtIS+gBxlpWJPXLb2wkMMk3qhHmXgs8qbMfZn6Fya0eRKVcxZZVT73rqnC9whGz
HUORKsYGFyZZnvwx4KZkhutoWw6wZoqGYg9NgDYJLhiq8nF4rEYytfEsrrivaiAe
yUENvsW75ufWywTVQyu54OVh1ZgxZ26GJXEKbZ4FbeLuuaVeRPvA6WFcWrjCiMnc
qUYRqTHHGV3ktKvJzLg9n+iBDNHRJQ1GlKf716EkmmlafWOLwE3OBf3BfvEEj1T7
/lbigs62tMx9PiLYUb4kdMk+7Kt7FWtVEJwVra5di3qOiZ8QlDFG16zn3cLIXHIW
JO+jtJtLIcnU3wkkRynB549vq9YG/pdYs1vds4DCPqtapw6Csm4H+MUV7Fegk9Bj
ezIAhTBpnS0CK69NaRY+2BpmyrJ91fM/xKXPXavCnPB10olO7lnD7DHlBScv055t
KB/RHUBgRfwzVCJlEu7kq7PWFwn6OgvdVbySLBlPi6a/7Yip+Kpbn9uGnDKRIKfB
znNMxOBJZ2RmaMjhzRJqVkBEEvPnDRIxjrQi9FjF1o32V0KyA2XVapPIBtwMRQMg
B95k651WiBxrAyGb+0ClHR+sRbKM1dnuGvU8EGrCFUCfzD5OZCY0bjNPqKeQ3Eby
uDMuEcdPt1IqZMdgXHVURXeDdob4cEXYq/yK9Ra2z0k85ancTlCux2jyAkhSELn6
zrNL7s1t9dZlWA5qogcJcZKUVTv6LkM5MBnXB6d38ULNKjD03pv0h0Bi5NXp3raR
jhn6atW3n25L5NivlBRJopQOnhPTYtfTMrpYbSxehBm/gcdGvgKkPbSnFUSCT3K2
VvIIpU8JmTLJ66woPJrfUPmUqyKhqPC6+/vdJ1kaeCNxLuZoQGaG3UuS+xpU5gbp
wk03UBhdipUxeo3C9QfC8FBo9kA1H6P4+0kQxnA51bX9rpMWJwgCPjXpABoPty93
+7l+knB3pRg6/RjLb3jNJCec5DjE8kld8tWgL0hgNEBcI6l/x7gxIjbADPoOyEFF
gsz+J0fPkmOEpoXkywBaxctlJ8FhCRwqIfoey0O4qRrZY1V+sm/ZEqJe3BPYO7ej
SbBKH7GrlzbA6gu/JURNXmU8sJtoAaVDPQTfbW/V5FZCMvFrq2UIZ2JOfxfB/X1x
FQY6M6PK4c2G4EmhEB8J9djFtekvPmFbyFdoyow0D8JFv1ayj3n9lS5rbND5tIp1
3hVu82ra98itKhHQs7hHENQPz5YjeqkN0wE+HpGCmMVX3yNHiSNmCcO0WXRoFNqI
UPMpayXsoHWIeW0JcKg5yvZ2tNYeQw0HwuthrpQGPXJ2prPcOllL8DvicCPS8rRx
+emvPfVYgfNWFhLqLek7TCeskbRvk6mKUTOTfeDickmwHq20LqxJqUCpbbVVqMvo
i7JZmyIDHVWFp9hLdfpeRsPLr9dOs2xJS3MH3XoFsmGB6/D6uFbP9RKXwjOenwgm
b6kcbXV/5hZxNanA2hkSKSFB6D2Wvuh6J/N6YjRZENH3hexpm1q2JDCEEh3ssCQv
+XHCPN0H+xYjChgUq37jweuSufyKRBTz8rH8S9DWvQhykUl40+0GZZeaARFsoFVg
2GieJ7sU/EpVhSPzlB6SG+9do27wWWPK/DL8PoHaqKcq2xdCPeVQQ3TI+CTZE/IK
7c30FHOkP68X19W0/1yaV4dL90MoxitkSEkjw9PqpD7QQB5QWd8X/aEDc7areUzH
qYp13aw3F91sx133t5kPdon8ZhkWtE6qaR21oG6k7lNVhGzMFz9DfvtqBqsKlMhY
rX/PxYvFLCjwARCYCiMp6SOpFeoWU6YfxphS0pk92qIbPxhahl1cTICPoOq7BoFQ
1TCcJuUI76IrIczbhQafm7YvqQmfFjxsSsdRuRHaxngitKf3sPz/lyjzTbJfm7HY
RHS0GrrHb7NAbKern77hBQufVKklzHOR8mE1hQA2ZBx8vdNnO6ORSwGIicMvpum0
meMHq3YjPj8FpFFgXCt98XU2XxGi+MuEul9iwMrdvkm0Lr7TkZyp3bUFW6Y5kapj
RaAcUnoC//hfhEpbNQT/Ru/dKTDRnEilL74FxBSi+X9yScd1NFuPUpzONH4tuLyZ
c9ysnRcKGTavXQ61iK2utWUqOnAQcSoDy0Rkmmh3sSqnJV/AZh4SZbPgi22/5zSF
LkZKUCx/+Dn5S60jFcKGlC7SVnlGVTmDAMFxA9qzht1LXuolwdcb7x5aPO+roVxe
NA4z4p4wkvDvVtsxZuE4iDYXh2K6bttlQCBtgExyHQA7zEWItszlHMPN2tdKYqtt
fmPF8Sr2qpsYHQNUqM5oM7MbgSIa+Vkf6juHrB5uKxWsdeijWv+2tN7vS5gLNgS7
fUOamd9fw9h4cPhgz88blk6FBtVGbZlUAfo77Fkj/h3KO1GCFqW0PUTTSyGIwXNm
/baG/naMTrzvTnnombM3LhPitXMvyg8rOo/L9wKJCpHUHM+2fChXkkIxSfsPPPyQ
JbT07Cxdyq8+/NOew7AmsY0cfPI3EM2Egs09QcVu++jfGAUQ/OF/mGDrPl0fABaq
SfdA+t207fsw5scj4HuHuRejK5rjXIvwApey3u4CltD81DpOSYCEodK+28lEIhQQ
jEeCKSY0CelBvdQP394y5jHK1m1T6T6UtzZkRt63jBDJQcdWjCFx6bhqFMhh4Hdg
Ej5hKrywEA09DUaV2Ht7+ImSs+yMc67F7leWNEPUonip3bM9cXjjFW0jUdIEBxlj
a2MpjPu+HJ/jxtHuuuR9lIAS01IEeRwdAyGYKuEWFRUI+2Q8vA+XD62MxA3njAzt
XTFnmV8fcBRzYIWZaZ2torO+NBBG+W9p9ordgIrJS5EN9/BwR7BzIGG4VlBbJDy3
dsgAks//tnC6M7wCtZFByXjpChDzNQg8reQM6b/jkNwawpirRgapX1xc9TEcXXyc
FmirB9WAV2epSSzljPdIK0M7f8/F/rZeoCZGK0Y2OguWS6oqqH1E/mMlNBlOL6qW
1r98QIWXpcsUuiNVgSAr2WG45yBMQMbtWLKry3epCKm0PQ5iSMCC54Lo6cvimtJl
bciHMRT6gTD73cuSeDL3CtdmI11gm/v5oOcYPIR+os8aKui2Or4J/sZJnIW9RL6j
qYu61NMX37ACDV6sLMa+4H7uwLcrNy5OH9Tl6nQAMYIoR7NM6cVuSVSdQ5erXrnP
j0pfm/pmTcUTves875a4Z8Mz8GtdWWDhRVaegS4axMCO/9KVVt8J/yzx+Yhly5cu
nNO91wXHzkFiirMLxsmSfXzXXYk97i5Mtahq1BwFiPSa4C6z+Gf37T7cBHa0KYu6
ntBb62OyzqZseqbXcnGmnuZr9eT82963d2Qc69bqd+oJQ6IQdnNKG1SwN0W7jEE8
nPFEkkpUlOCJSqC5VXCwpgUyMUYqBpbJN4Q9EKdzX46uCRYJRNVs4OYI9pyAFLrv
gKhlRU9MI3xrnBwbkiXzYd/e+mouBw+FNzoM6IMRBrCRVw60PfNlAG5FV5wc8toW
vEWZGuiSBoPCyCDOd38JPtdL++XNpJkgXWxFcgvqfDq3OO4zKJAeSNhWkKyGYsRK
KAlO7/GujfLO6f8me2urmsZgi+GwlS1m6CKuIxEeBqWrqROnZ7n3n4+k4Ye5wXoK
MWP8AjsVmRWYNkYscIlhNleDgETb+H833zLTaDdsW55137xx1MHAfAy6jKD7A2k6
JrhEG/HBvAT4d0YGYxz2Rdo7Le9npv++b6Ktk9hR7oJE6mnxbvoAGS3Y66RSQNfJ
j6nZXC6V/DfHnQvDYBdN3woC7wKMMVz4l+loz082Rd/qdXkX658Q/YEhu6AXMdVW
YJkqfrymmwzUWPpU2j4dax7DTwOJkANKgnvqgkwkB9e2hAles46Sx0S2pkylOF6W
E6d+QV7NMbGnxdcJwI906IpkGPcziNB/9936f/NHEGpakaX2hYXSTxkD1BztE2Gj
mnscTmPgIXUgr/aBqn1IyOCKS1X5+A0tcPDobE5t4xoZX7gVFF3M8dFQ2090796H
lfVXRRLTXd4xyx2j0V2D+03qN7CVNityPQ7u6c7LWuuXd1XlGac89ZzzMGTDea6Q
f/UzGk1F8QXa9XQdWXBlptExdZ2KjOeTbWhFpwKH7w8Zso8aa+R2aCFSxWXpd6HD
KsD3v6IB8hpxoCOWGruGelE+6z8fhR72Yy1CxKrD1RKdydGBgpRjJ5W6yhYhrzu/
hjD5HMRP2R3nnjmiOjAlHGHH395Im6Npi8tkqVPaC8BvWlVoLSqd11jfYO5AEGEo
DiwiHBOJ5KWCtlH6T6oog60M0u10zTxML5NCnH/kP6DZF5jQ+wRres5jRzRp/NSe
MUkIjmYshzPLJcfCbYpk2IGeIpp50e7cOkqh9Je4f1412o1PnrqNO/nJE/QWb8ws
6ySIw8F7tAzw98iDla9Dk/TBqM+W8T3GX/zOUwPdUw7gu0FmNqko1GAIr3avnyU1
UdBGgOP3gNenyaGZYLFw4meLZ5xKjy79fwmKrtsVgXvq070QkJspgiSKF/CS4ZeF
WEuJ5IPoIHlC7k1DPqAtJdEfbK5IdBomdR1/xE5KgBukETwyFNX7rkjNOZn1HI1f
bPsXMMyWjJQag606vMjwdfvavALwEhNgS3n0B+B6/q7Wxdko1vYtPhnZ0xTDx7m4
LDzLMXB7pR2dy2go+nDfgOxhDbRbkT+5rK817h7v2l26vZHvpruWAwPBpMolPn6J
0wI73b3I9k6/8vvKAP9kLybwHPubiJYD1/bWiC3jr+NBN0gbW1lh3pcPnMxAYLGk
KLpi0OzNAg3P3tDMQZbzoD4lulwMUetVxj7RXzn0GgiLi5FpZhseDEY5Nq6v+/Jr
M/07zi2mzBNwne+A3rHSX8wl0Siiu/je6Yx1Htfru6B4Pwf8x6sQuCYeo1NayiWW
Kgu2500XqdRCo3t1+yj8ZndVHi5q3v7IC+O1IAab8+dy787K2BRCOcmbA3v20EOy
fONTzm6uWYSAhKJvplTn7IxrOE8W3NCrfXKZ0XUW7Q+sAHUFy9KoydJzhfZqAtkU
PysD7i+ep9/j+cVDkp/HrNraEJOjKTEhegGruPBsRsRnmOvDsSMTuTD/ULLBz+Ug
h1j7jX0bY54vPeXM3iHZ+uFkYS6UN+YuqEctAc7oA14eECz8CjkqlPeQDESmmtw3
7ZToUu9R9RCHkXXtBn3GAOGI4uye0gBjYFF7mXioX4L3gdP3e832GYbI9Dy8+WKV
PZP2DO0ah57ezO2Btkj/HPZP5Auc5roIWyRdoXhYbFMpHFTF1IMa3dQ18ZUu1LfQ
hhufEtL7SSM6ntDv5yCHDd9yVdHUKT4MkE4m68PMddZsPjozV95pfru2gEvkEAZM
OLYUsp2/C7fip5jq9XcljJNRBGPIhnWWVu2IT1FChnoY/kDgekvrOFJPuhG3whGm
TycgY4IMQyEn5IPYB7nff7NGlwFnKN3dip98n4qZ7WeNn2TcO6tnaIHYmmvv989X
zh+3l18m5CfI6KBFBjtqOXeKjrpq7TCQr0qzaLDO3E/c5igf6E7wa7iXDlgqwA1b
guHOC/uFLdjU0m4bWArc7lRFszoDz01MJamxEwbEeP7b1YHidqPS39te4yJzpBhW
BjzxecJf7sL5+OBft0wN41a7n0Sm41r3YC104GD+9t2oqaBHvkYiBWP/5CKZY1qg
aNfzoEkilw25myXFkx/U0po2TxkSVFN8tnLdy6phH2SBUth2/l9YISFAJAHH4WYV
OH/01pZPvqM4FALR5zVs6lhaJdHSgWkF/px/QF9IjfVCZAJ5QpjfSurzakpVHjGE
tABuCSZOOj1RGdy6VKph24B+IsfOxWgFSfNBWMymACbT3tfpkG6ReGtdmQDHYZw0
gavDmM8CNp4NE9CHKK61zABA0SKBBowhV+Ba1ncByNEoxAh9Y/s8Kx2dcGON9drw
UcICkSSapP6cuYUunr4fw5jZ6PuXAfK17LjjE9kjgEMZ8yy4gn70Zl0e+mo6EUgf
WI1lAbhoVXKned6BaLz0F1XVd9s3C+WJt6cStbDHmhllwWipD0YaL4x5dkUH5paD
ZadNBhCagyklcghKdmTlscDOGaGj6eGnluOU/eaui2s/Qu1J5fyc0i20H/Gjulnp
Fc7ad4X6MnwywITEYvv3boma2T/0KrzruvL1xitCENSv7R5lb3RMTHueYsHRSEFD
hpiP94quBTg98s52kQNvUeX5mCZmcllWZHSDUw0t3orUUMts8uFwxlfm/Q7G5Lek
VwdknWpo1j1Tu0olPKhCCyV+/+3JaRdJ/uHoSRZNRX9jyAWnnpogWuYXP7h83Uvn
EaBoRMGiEIcP2NFOn9j/2MzGLkx/M5Ez/60zs0H3PUeZFqIjbjBbfN/9cbsuRZn8
CLcBs3dWE45Z4RRtb3mXCUkHRSwIhQlofuxLdK4onyon+FdL7Am0iGQ/K8Jk0771
xDJSrX3vN/i9fStxRNLCZociLQvVBNYcT5RYzbzppcG5EyqisRa8l2DB6PKyQ7Dz
LUsR3skuOtlCZhDJD3E7uCd7A1132nouvWS9u/8esAz/SR9H0Lp39EXk/P+YKGvv
R/YQohDIgJ7/w3F5cAM4Ulm7CTMi77LNXTSzznqqFW1A7eO1sxUd6aFtiSE2kfIq
ZQHs909yPTlVI/Uxz5HP1GVbeItEqsuQDERurdeZwg0E5uQSd5Qr8RiEog8CwgLY
k/H7EH1Obj4DKR31MgdSHCaMetFsnafeDvvT30P+4KCTlcO0aIBvqFlnLQ4vRsVo
0QmDsNhYXWBSjcPnlTN/8yEV3wv55IoE5eMQDjzsK4dqRI7VG4w532IGcguMe103
2wrqhDqvT+4tYcZgxdzeJN/6xzEkShPyNxEOXNox/pqfzLy2zIk8koEpXPN1jbJb
4/OIdXc2ObXi8p4i2biHOyHHkbrUMvbe4iGUr3tQb5Gtip84ivhTn5KMDQ4yxrJk
D+szRq6lAXZurFAzMwzJ+0AjerDVo6139VgVKLg4CBzSiMGUP+kSDMzFQ4oAZvoF
kKvvpx7GMejRv47A4h7osSfKv7F9kX7bxyzngCsmgRROsZq47NbaT3RM9TyFqnGM
1YBs6eBzLCv3n/1tDMTRitXkIg+wLv1Q+0kcV8NfKHD/CT7K3eClllKrNgEmz1zb
DYpXWqnY4TIkMiiohPlOSrOZmCltc/7jvZuaYwDaViyYZlLMIJd1CAThtyXZkQlE
P06Mit67vW2Su0KUXweqKz+xCrATgqzuDjypTvT6HZ4NJj15i7LOxWSsRH0XdGYy
HGc2X3AKtlCv8MkBa2UyzBwEta2JVs5UV9Zz4AT/fvLLNguzcQBEhcj8O+nUa8jv
3kRnTQigcuBUDRv6hc7Y6QEjfCpVqRbNT9Jc7kwG6vvtYpWjrUSZ/ese68gZKPcn
X0jf1pRs5HfrjuPNYkHObBAaK0UzyzWOdGkuKGspFbr7vlugngCwY8PLovJR63SE
BMYQVQtHuSSt5RHTKLJkEbRnArsPz5sqc+dky7Z8xB3YDfiTohUSMeFohYza1qws
1kDkLL1SU5/qlnuBSCaU0vZNeBn7uJBRZ73gLi3iBte0UkP7aoZAib9TfNKmhkJz
8BxV3/Dixu5DtkNZQBG7v7JgMvtPictG1HBzXkCh3WHe1TlyZIdr1N1L+NdV8hzo
2oZHXdndVWgpwjgPROAutcvqy968loXxHw0Cp/vXEVYfDWCEP3BYiVYccgt1axS9
3CxVEKfO2PxaAdE/vUWLxryDx94IsNDxUDXKWUDyqrFTtMqk/SaPiPQr9UpfO4Nu
ULZe+gIdlFyDox/I95c65oJ7OjJEE+yADdAh05ywCoZFi5XWQVxbclr96y73XaYS
xvbxYJq6iEepujsOBfJQv1agovCLrIjfbGXkWp19UbSRSxuomtSjAxna+pzEzKM6
ghhk7yX6XfRCzMOPZe8pcxSwkVBliOm5+fOH6MfErxUCEOM+NFx/tMoG/yM7kXzc
shjgixl9mArk1ahXcgCwzY/ieK9iR3rrzDfzU8UY9/HtSkT1ksxit4gGqGHd1X5g
mj/c2A3ZVuZBQ45dejtfq5lJ6VUEEXH4w9PZcvctFBdVuQLJiK0PuTSHzawdap4s
J2fvNedxyem6YRpvuFg6z3P4Ge9MyLNeoLQSNsF5niFSikCVs7tuONEHWakBQKAA
pPRyHHwCOI2JrreUNJ8c8NOioHeBRwB7XHXDzbYrXfSv2Rmkf++JBxHYuWrx1Is2
BODQWbPRr3L7+rNtuARsFrOn6Rxt3DojMExXfv3YJZCEf+DUNgGGAimHS07r428D
Kn+rx97fV2+3Ag97rxNZv7frpgqYELQ4xyuyOf7vFAxFHChJUsXqoZ0UqpwW2oE2
G1H6pHos4aLhkTYzPAsX2RT8l+h3ZC64zsMWTkmoaeOO1K+nNoRQEocWSxaSfSmN
4cv9ZYqTKuKbdeVO0GvoXoC6OXsGtg8Fxb1N+awRBbQNffVW2lV+4k8vnaqBdMa2
8vZhpysk2KGfIz565ZTLLG66k65w0a5ocELmHqGxVgm27qnDf0EksXe6RdNrgnDI
ylK+pBEk7PDiw/bwBJ0B59JWdbYhbSXH/9mhENmvl+EkIclD67wY64tTcPUt5xVB
DVpQ9+GH6akHOnVu0g2VHIqBVKr1Lfv2EKU2pnhJ51vcm8c60DpvTpj6GC3gb4NO
VoT0K2YnIbARrU2jo82K8bQwYIl4sblAC9uDQ7UfGASLWhBR2oR1/uMs/vLIp5Qh
onZRdHzRD6CNdcb/Q2CcKEMLddJ8vpTiFonMMM6yFfvPAVaER4zksiSDia1/Hct6
JV8jh17l+dFh+MAWoCPQHeunYOz//qdyZrNfXKZPawHNRpjy1jVG/3SjjAW1J1Ic
ssdPkHBWKrmIecMNRbYPyHlWM2ZZX8DTfTMc4e664DLzmKXeJzCeFoG1ojB/5egx
iMvrf3a49JTl6uHIx1/uotPR9TVEYZCHiedp1Kp1y8dr4WUjmwdna17u6iz0UHyy
tDKg+5VldaV+xGVzNDUIGjpYZIN/IvOU9MhWxhtmchqmc1allLHyCC8xSvoP4i48
TFYpHhRaSz1qJcoxxMe874U4dXKNYVKMLcHSvEkcTvHmpOpkaYsUaU/xqWhqDkTN
/2uM+B89jRGw3nEZYsF1DqI6bvpnYLZhqirmzaUh4o2Yojqzt8tA9HmIgSj9gtxj
W2VGh5OUrVHr3B4Vp6CPJS2JOWAumshz7TNdmOTwvhlu7vgibgld8xVBMhPgZISo
58Y26YLZRVci1MKWvvPOG2NahoTl3O7aqYja1a1ct4gCyL/R3gbk4jH3rmOzYFnE
18+GcgG53mR9CXxXWCq0zyil6ZZO+X/6a3ZTwPkGc/WkZhrRkAFf3tQrRwC6ecm9
sVDm+VkmMysqBnvsFndZo4+7ql1rtVs21aToyUexwdsB0295yp4uvI1D+sUoePEx
w88M3fLkIGNFeGVYXmEUQowjEq+jzcHnjJJ/AnKlFCTVZK7CgUSGU5oya7eesPhm
keED15ymlnxaC/PypvbuDKpg8RIw9uQxZ87G9SYOGbs1A5Oc9PqXjgTKp8GSC1nk
S2LrgqF7cFuXfQdrUw0uy8cQDm8Zxs1/S/WooJSshEalHmeY+gNgVeZ/mxBlA3M1
m01mZvKi7nLNjbQDMeL7XuJpkxEDPr2XFpY9tyYiN87hFAIoruryMn+89Rta+1Gc
ThBo32eI5ljERYBBZ5K4lpPKVi1q7aGQTXa8CewJIoWbymtLTdMVuWKw2kx3GRef
aPTSu91UKjgNcGXxwa1FYZOXXGWXQ9OUCxaanmC+OQ5BhlMHLroqS5qYwL9dqymx
uFQNrWwVNqj0lE47ym9YabLBsz7WeCYPjOqxAbGaJjRjChxRzmfToDh69srdkdea
GUkNXaDjXIZ0whKC13ffkl2M6gETWryf75Gm46/6Yj9RIEeXbxSQOG5KWThNXB0W
rSd2UY+InalQiK+HYC1U2teRlAQyqxEwjxMctN31lF8Cp43cKWwHTrOOrSPMWWDe
QTFohTskwR7huxwQJtyR+DxClIIH8+62dHYMsrMnQl+TsH5pfo4N87lU5E5XFiVF
0+4XsIDdp/kqvOMc2koNqB22/z0eINb2kVuKE36Ut3xLTdb2suV4KaMZv4AxhNqh
HxEYg1n8zZnNLpUjCZu6SR+jloJeoMSU7J3whH01VhBgkLrVCrt7w3wKbLlnpzdM
sbnNIClmQtwAEVnz6UNKjChNlqzI/kgRC7jfN1Iuitsf6rhXSEuJ2HR+JyZnc/B1
Kbn4W9zr+NB24r3HvvG36dPrZ0HZdC6tvzHNfT+nETBFZ7iDNyoa+Il1EwdhzdYF
yc6ihngFdr/BnwTCbk6ds+GkfjaxGRhNhHERMpHbC4c4v2Nd3I1zKeXlcT8WyzvN
JHaFYAWXUr3XAqJuEpCxPpwEmk5rIMZpdOzm/AlquZITvI3p+A7BwLfCHWqiGwLi
8IIQV5dF9zrD350bDtik87J48HKmKPs8WnTVytIIQq+oJHOl+A3ss6I4NIMXEUCA
UEPAGeWB3+LNv1QPg7UC0xzBYQtGChYlA6Bf8yubtwyYjD6eHNS/lcksFzUQ1QjC
3XFp3szhcL8CemCL1cDACyYRT/P56y/m8f7TRvqqun6jAgE31qKHUgkFLr1ltNRW
pMZKR/64r9eHuQMmojL3pSK4TG9ChW9s/jqp3ubLnxfjxhrgU+CsANgO/gJ3cG2d
DqSOCbu8nF0KPpr2We+FybyktmojESAV6LmSoZ5k1od9/yhXSz8TldR822L9nHrc
z4PxcCWzUip1YlaCHaAYZIbmQdipwsSYQMb4wz2DcuZDQRG8h/hyk887MVBuiL3I
ayxxujBqysKotGHy/2bqdHeZ/K/9IkwJ6WT+TKwUpV0MXGnxmdyAYhAmgro8wUGn
iUqk8H3l/LLkTL1DD67CtLyd43kRQc9KAQx11QJI+dzpvkctepL1pmUV420XZwLp
ZRJ1QCnzMtrYDGZh8VHtt7jwai+6Mztxs4+2CC6H+vQ6WBcmX2DkIal0kTnExTJa
2umP6ke15qD7R7Az9T6P+EjjgjMlGdjwpDU/chjWJztuvIdtWe3FN4S6e/K+3m2E
1OZMDQOdRg+0wGs1uwNNw30Jy8Oz5zcWB96DPZgtQKZFRwvuZL2fwtZmY0pGC7SF
ZO0B62Hp+xqO2sv1R6OZkHUXddtgkfQ1MQh26Jc/i9cA5bcKeWu7/41thRCjdbCN
LPQHaM+HviQcaGUkW3zn+LE3+u/LxG1SE+wt+bInydjMI3iVByjqbOAu+ilkj7aS
ldztf3E/mrOx9GLDCHk6ALuQubv88kUwQnwditR9Ueli17szELUAuBgDUtVnVtC1
OoaKzwxK36IYWnsGWf1RE9j0btx5Fevv+EGAzwQf9/6Vt9H+TJSqsL2Ly3I+cya4
hBRble2vv6bkuxIgpda3iT9gu+DMwBw5wABnIPByCSFiJWUke+ILnLw2kd3Vlt+p
tW06YP1HzWbGwHG+oGifB81X85JQt1JPZ0zIWCNIqbhIY/i6bmhV2Qtt/TJDeHqB
zLvFjGw168VnMksz70Bqlqifqu2gsYSmH0XcpT6lmDLQR/DiCFCN3WFYJVUu8VWc
2uhglOuDsPO1D4bNOZrg7BWeAy8s2I3RnF5i4+Un7k64GhDf3mV7bn3SMEbFMVxs
XcsLyZ5D6YJh1Jsrp9KvyKG6bLAGHxOmtMjE5BN9xYZNwbpUZhF2KW4Y+URevOhA
N+iG6bjuv4pci399zLyesul9Xi42YXi7pXbO1SwJzhrIa7BNqiA68uy3LtBHShqh
/UY07jHC23LsKhVlUevc/+nnN6n3rct2rSupuuWNRy9pSkC0QA1Bh6X+tW+SBB28
rjkVVAs96sqnCUGA6Um3hvU1gxpNTokTci9j/ZHz9ZAB9zIgjI8r17OWKe++KExR
PK0tGKJyN62mqZOFqDnURfhxK1qUOXyHULY/jK1ZfhXjj2bGqdJF+jTTcdtep9/t
VX+Kl5oCa0Da7TK1w+wYrU2XuF0eZz+hGRGPPAJawEmFMRTDz5muEFe6IxLyFsup
ZqnRacVrQydtTbcA2mu02glhcGul7BATYoEpvazMspyirthnN9HqrPMlU9qtIe4q
Yyz/Ay9XH/FSGbfJqCwVKlSDac5SOaYSYEBlVay+sywKtp2n49qpecLt7OB0oT5j
ZTyUwzQkjkgZP0NN3CxWDq30NvtvIIg2U6yCCOB3mDNxnkHTRqY0HpN5sYTAouDt
r+1TbgEdfTh+x4cPjx59N/2D5Kch0S9T7d6/BymBsHosBKsrje2vJm6Qb2Xq6jIm
GlmMtc/aDfEmxco9tJ4j3e/Lj405i6GU8V6JIsqPohtzN3JUT0r1SyCpYe0YDFQY
3Epwssz8euZ6xFhQEMrpbt8wVjl4Oz6cAlS+x8J6RB6NcpVO0gEnCylZgiLHzq2q
aP52p8FaRYc0JINhtEIsikzPCjtV1Wl7/yyGLjwGCyTzEyPDICWe3/C2RrZl929Y
/h/27Rptj6MN3gYUzamvCnv35FXGLUP2vCFkh/g4OBXfKAn3OhWJft0uG/FMyBcN
kcB9bvOUYIJlCdX5rLUQkDKfQiHmYRWbveXLxrlD2s9OII1caRf6RU7mcYIwULvZ
XKjjQ6CjZPp/CW/1G8X/m7LgbJ8wU9MDMnfBbNyhGpCmAieiaepngs6l9tvBmnJ3
RHAPuptuZUMCDyuKYtI9mN+vY/+xfnLPOB5kh57t2bnXkkryjsGhNUXm4tD9eNmS
cgZd+Zj6xGwhJPiA72wNPRRywKcjg7JDhOQTPVv5X2Ffb6VX1vJha9jAA5ix3z31
7tWgiv972moz6sPYaxf3p0cKhjGFsRcPEAG62Mjr6efGXcAKyUDUCpQ05oWOf0tp
FI78yRsciyhu7rl8kahjh0ufP+LIoLHcMom45DR85foZviYNElGvB8um5U0NKZ0+
dL/kfpD5EJUqCxF7bihk0gmxx0uM4iIzy4eQnRWKv1t5FszQ8w/2C/8pyL1apQPK
0Idh63d4FIofqAvUvObLeTNRD8lNIzpTxhzluam28OfHnsOOdj7UDB2ub6L+HxbC
vA2ezUjNUB2qunHIgv2znwjtlpRkhgPGkYN/0WbZGpl+0EMn7poTB3OvG27GTSUs
Qxfz0TmXFlsEsgdGx+k9GCw/QhkPwdTJoKnj6s0YWHqF3Eu2ZA36gmi+D8kentUp
B+hHMGSw8fRF+N6gVV29kUWlJBTUoZfmVu1SfKmxvIjVbyhkyQDNcr2K6p9F1kwb
5ecFD24LiTpGQ3I/n9gZAuVAR7Uw+82QFUd9RxZJAX3HBtnGc97WQSo5pezSus3L
+BDa6ruDOLeQ2rzIag9TounGfd9g51NGFwPcUo9mcKro3tM/LgvCT9cWPrsYxMZs
u8ndprpYsXro19vH5ziWBd7UbxvPcanEv4zk47/6StkQDeasUQ+x0CfaTeREwc8U
3UZIpBDExLYUkvTuAJQhAS+eFz4sjkYjb4vNzfihdr+mYoDnxd9NVuiY5OUxzW08
JdFix/uGiFzjFDoxbULX79LbZJKXoTMSQIE8piHFuUW/DAmTQ5jPfz9/EvjDTRtQ
KtVnQCa8Qgr531VZJ+eu6pRAjWa3W4rCBtmHGGbROy8+Y8p/7kFP7C3IjsZa0J7A
/gFwA0KM2LSWymtv2D+szpx5tqSmnY+GItbmScNPMA+cYnSJuxmVGynimQQQdXJe
/zpP4Vn04Gna6ChNev2kOAGHlWwt0H7WJROM8+/GtAsVzEGZnfPdzxvklOjMs4oe
1HRngw55qGOU2EU1E4+V8VdWADFcRss/HhRcl/VH5IZ7AomRrLqXyTRyy5kuKjqk
a1Un3q8uKZLI4YfCvMjX/J9CRvVtiAtDqQ0Vcfwya/43FwkgSVy2QYNpFH1bBidY
D2JpNqh/M9xY4u95U0A9z2TU24B/VZcbzkY4qVVrfJB0/AEFs83dxAP/yWGbElId
T5YzlhlxfGV91Bz8tbw/uWKKYLUjcsZPP7fMe+9fIW76WqW9SX1ENSBmzvL7tVYb
UFHFpAEzKcnUO4dlXv02U/pfxu+SvfhoK2OnanJSAF8mlCBbnmgRkRH3ldhY9tPH
oYxaYx+qQ5DdHrFcHw64PjxXfVyJ/ityA1zyYZVgSeJHGFo7FZpjInQY5L7BB59t
VByePHyGcWkfVOn+iOY19ebVe3Vqm83U8uc3dqO2PqI1URDvRfJCdg3OZIkv5uJ2
Lcl+m6UY2ehRgaV7QXJKN3AFRJwJySScJpRwQFgI5/C5q6pDqUCdej6T70i3u+2A
FrIpmNcyUcT43JmxlmqJ0iMdFESRB363EVgUd/l6H5R5+8JrK0N32MhiBb/TK7kr
B9h4s7sSvCX7Vk9Wz6IgzJuzcc1HuhX2zBbRoQlDMQaiR4Of6n86YpvorZcN3UF5
AWqfV5vRQtyjGkHh1z6mJLIP8uRQhpzScvIiBwXNldJhGkeL2AqIWslmO57oqlvk
cueCgMeoD9Q0i3WPYz768+5qdbg0ppIQbfc1Cm/DU1VimzIQl1xtd7+4Ms4fVVX6
pZRy0zOB1R0th8oj7nDLWDuUaCujIZL+qPTGVfRpEsytLDzLz/UpDFIpeylTIhKW
IPGQmswnUhEX7cRepqfA8KECUEqLecj9l8WilJ45tjm6xzdbCUlEfItNzkPE7BBZ
Aq4d0/QtY2kXhLmFl3zugQtevwSzr+vYodVY24Q4dSNLSGwMXE1QoOTkiIYTv132
6WE88qToMlvoQn0uY3ar2+O6Fy0vYtrhDW6RQj8QgiY7IhUkwUVjcYDZqWO9wiQg
rZb1LS2M4U+hZiXFW63tDUM4pdxKjC3UqhQfIMaBlJBtQGbRQqwQlP0sajK2jh4h
SoHAAHFZ7tYtFEHV7qR9CEelLuIVf5U4/NgzXfMcxEQCBpRKgWj+12t5cQzfe//o
+CVQyFUZdJ8uwYBX6hBZ0QwDlG61Vb96szF8FHrTcHE+V+/htf/Q2OJmq78DQ42x
vpuWUzdtZaVxOE3pr+t6cCVWiheF/vpBPgwkybx6IQuYDbEINW6A3x2FL30by3Aw
adJgUwBXJ1Ce0kzmyaMq9VEB5cKVOMr92rPB97QYQK43NMKzzHlz5VA1B7NqSgv0
16Mrq9mh5eJP4jd/H/9pYufvuh0udQ8z3fae1Jf8O1xxmY9GVjiX8BVEAyY3oIb8
un8TwbuCNzYRGizJuBAV776ZONkJAKa/mOoHXEQTkptvJztiwz5QeXwFQi1AgDzO
GhPG5LpYipDsxh4BWfTwn84Opsj0uB0SWd7F71y4s5KnmSGStgRukUzA1Dn66Ppg
Fs5XLF/Wtf+ZCf8onvp2JB8hJ6yDIz4JDsjwtRhNIxONElkVrV96ajPoylDMuT9u
NMSgDUSzQZtXiwUBc3m56RNapuHnSgEgrlVM5ulm/sZAgrpvTMgXVjo9ErkLE1ib
E/yZa5llwpNayvFbICqPeHin/rKf045lusmRayISjK7eCS0FjOr8NVmqsTG5Q5LU
rQecFinA088P4+5eKDW1utXbCfDOXC/2k0IQHfJOWgCqyPdp6Hcvz7jdJkzpQ8U8
BIR5jPaU+ZQ7CU8Z8C+zqTFDX/pr4qrTWhfkUvob/1aJ2m6wy1gYFigzZOWlgGvQ
fSvKEy3HPaJmqERzmlXYktgkRZajaBi3hnuLNlUiY0ibiMt1M/bWDH8Y6M+C7mfU
Dxdd7ypLdQ6HfF5pX45sKPvA4B9q45mfhFrZIpCWOLLH8GIOGPZADXfF0iMVqiY7
1xzWKfy9k62SED1g0TxqN1mfyTSnTwGHZmj6NYkaox6tqpkz41U6ys5Zf+487RZb
h7SAleimyLefs5vfQFBu3pp1GtmJAWm4RQuK6RkzoVY7zshjUhywyFGbijtmNz1s
jdix1a9QBDYquPThWlp32XE/UBlo2v/8armQjQI1HOOuX5ziJzilHaz88WHpBS9Q
ZQMQVXW76abWD19xZl+jL2XOrwH+G5cAb/3wdRSNL/vz0D/Ed2s/DlvKRgeG3XQ1
AqzC+vTyFqNnxmsUrDTpMBjJ2a2X7GMBBsjYps8uekZ4r961d03QbXz2ydMbJxkk
LEw6prh8X2CidyvyD7CYkCBnUPEbHH8rJiHuyN1oHjWdhkDQRXAkDfP0eTdXwUA3
SQ+mPMiim7uTh1TklPNCgXAtsviJmBJW0aZLUf9Ri1iG25jnLCYdaf/3dFZl1PMu
Hkz4rMpc+8EZl4fg9vn9qxBkMIzRid8NfEOner5io1oDNo1sl6IfLd/T362kpD2Z
tYzE9Avu3mEBhHsWpjv3+ql6tlpmWXzT6s56A1sG9xDMPz0DRG37xxsCjTnSTUuq
0jVHdUnSM/Ou6LTRu6ZD8pjQc1V46Bat4V1IRYVRlvpCRZMfNg7qJoK+WcoUERR1
LQ34165ktxx42oUVp0lmZ2HWqkx3eI7caqfIbA9mqtgV5W7BM0wGsMBpm3Iglgeq
tCloHK6N2ZmvIxhMZBewS/pWAx4DxWBrVVE4yvcs0vU6lvEQaB/Z2HBajonlGIvX
Flnb+LsdZmfQmbm968Y4KG5MUJnB8TPhHA4qlvS80rYAgERvZNh6uhyoQ+4tWmoC
+vKQJ98Rw4jGJR8YwnRCaby3Q1c2T31En1PnJTMbfWzaQ9pGs6s5P9lIsGm07OLi
weBXRVE2kJkgH1qXVtPVBuhyE6kQ4XkLxnA/i3wnq+3De0j46bC4FBdAhS4kn+GM
1XYi5xvtnLsWcZQAJeZ5EG5H8wUNw3gOuteT1xyqMb1OdhSEW6QRAf/TNKi9G+7h
fHblqPQa/bp7iII73gmJA05iUXkqkZGJD7q6I8lrhPUK10mVx5ZDWeYEbqzqmcjB
IDAEMkPLlgJxa8Y4iLtSlsdEs7dF/Y3OBxV11jnRf5raoOkcGWHScn/S6XrR0CoF
vwD9ffUhxYGNmeg6+TRyGucefa7keToyYkaFrGhP5d9reKno5fxp0Zt+DLniMw9L
GPH6qBp2tqGhFiVw9hyUXJIZXKgGE6vOIVP4nJFNv8V8c9C7fnG8X9xzAICxMcBZ
uoEfrUiY7/kACZ1DFuRUUzbsFCtHhhzxucYX+yvEIb10UYC83s7zov87d/Ns4hIT
M7MS7oS1EMcWSJT/pX8kG6WYH+TucOBDwx5vRBmb5GNmfQUqc6UNTDQKMk1epwLc
t8kypDkDzXAGfxPtWmQ78BXy8zprLNvEYtnLuAoPyZl/voqFmz5OeKsAYhkXSN/v
8hKL7Yd1fOfNYPSUAqn8yYOtTdWeL65ZFQussNc+xiRKGLx6LDNEnva1NImqtUsP
fGf8j+AUG2pad9f6/Ed/rhstl3XW1eQ471b+ah7uzRBuNyo7owaWk/qE6nXp01O5
AZk7kNl5+E6Dxcdce3Mz2y7kc+I5b75pUKeLqQbrQdOYsA1cahrAmKS8F5A7SnaW
Ssw5FyQaWtIZt2jXXeBWrGHLX+bYazuOyP0bW3vcP/xK4xhO2IHTi+xo4yyYTUBU
1Bxja5lGOXJZ0Wm8y/ccEZGc0m4MFvN45W4U/ixiouAwR6uOgQd8VOMo7PHm8mRj
yhRga28ryEIWILrdGdMnV88uDo6e6Q9S96IFoHTSx2wwmS2Gij1F/cX6esj2DvvK
kjMgL36cf57vuz+5RNrsPbM1PizD6lzF+QQRTW+QmfV9xC9k8VD5QHL4awq6pgfU
NxVRp6fkTEVVH7tV/aYkk7yrRUZ8Udkcap6mPRqXNkepC2rjeP3c+bk4HvwJO2ZC
dQP+7IqA/f3uSylVTQscPLWUIKGhtuaQx/ytefo2XJkTkj6NNVlSCvKMgpV6ocsH
LQGb/U48+N741UIrPukx3br7Ta5LTGCDQPs5ZKl6mHAEoa8MevirY4cWo80/ZiZC
R7xbktww0ldL80nXBHuGS865U78LMHTI9n7ijuaOIewcmw6DLZVgzr8ahXRBHiZZ
JNDeapYhZQvUNBpZI4YbYT7ew7ho26XSQkjsvWRhU4JsQdI4PiIKCt3xYsz/QuJz
YRs3S517cVp3xfbitqWqCN6lBmEsjC+NPGa6FIVtWR85HGHcRpWafnesmGItWNO5
E7JdHdJTb6rZPyK594f4KNbQfgCi+iiza0SntuCpeDWREIWCYsbsZv7J56upovH1
Zr/uFdxRMLWZlveOvXfx0ZMenCIqqrdrrUJC/LlYXrQqLs6HW2fik/QBUPnACOWb
aEZ2hN+0ejXXZ//8EIN4zALpQJslR10yEpHZAD//F7sKl4QwZC4YLFiaglWpW+Tf
K2GG4OSKl+WQ7NmAEStKqXm7FIbVo2gUKVZNR6YYDUTYrwfi6UvRrv8jKbhHWLYN
SIFNIJw18/q3l2YkXcGknnwKOT+Cewxkfj4gD/TyrQNnbDswYtY+mHMRSPvv29mf
mSpzub6h8qLZzpV49DI0Sxd3aI9FUlkbVneB0M3AnNrjwQJqf+DKnYLMLmdXqINg
3pfvN3z3Cg/dNi9D7YqpaOQ27k8Wj5LyG0phGWkhPldFJD1ULAOGgrgd0RlI6Ch1
Vroy6WUwIX1p9ikH7+/iQDUlj9a/D16FaNHyA6Aelhlq7mNUiQaNW9kujBcjPwRd
n7hx844UsT0bXzf9+zKk6KhYEO2JEHXvHtTLRxs99NcpKAhQ/rAgV9JuH4xPKpuU
Qfm7h3HX54YDuKFjLAmc5V85rHg1fn4tafRlSOKUzrFLA0yNjJZhLykEY6ig8dQE
C9uFpt9dDQBkZUWPdydWYgbAhXN4yiVzPsoW/nrnqSmBu7Z5T4E0auuBjjdDg6g6
nc/xClAldkHDSBuVennyzLQyo4/iXEV/yk6AaaM/yOXCQ4AOdcGoazMh5Pu25Llk
OHLOGIS5zR5L6NEFaql7kDvY1vNfWxQWzm6+XBKgeMZM+e+ZvbsKwqBvUq+rwe1P
RIQgQ3RgchVlv7VuyF++HP7RMTUWcvcnSWDxG7iK+r5XTOuKWCuiSZYIqINiAS+E
4UFjRPTmq8uUAb1hOZ/ZUFHIFLYZdhQtdjVDi/apDPEYnt0byYbLNoW5mYKD3Jtq
yi1113eqXXGqG0v70DNsmZLRSC54G3dyU0pJ8KeT5USy48j5dwSXk1kP9FoG9v93
ImPND5yvF53UhLGFk04zHT8k3k46ffVGvv2CeOxNL5N0wQU4b+wE9DX1hK8x0TJ3
X3VBsXJ0+/FW9smHVk7cpViXHhPaYVq+2FA7CgO5vyM2TK5udCN/L+vdb/M0IidN
yKz1YWCYzNk992+JHI9Z/ROWCv4hA+5kBYtgTXQtvG+jToyftwXKeA2H4c8EhOjZ
6mDYp+FU4OQwFwMUIfIYqBkdo5RVgs6vnapD2JtOlvKAyteCnC3RQIwNjumVAsL6
MVFxfAPcltFptGfaDRlyKErDbG8GYemPZqjR5no4VwHp6p/Avw4ok1lFBX/1InsR
r1IpJYBLKPyX9xgYj6+3QxYpsxp6hdGHSjJm69bBTeXb5JemGl5/vrGK7VCC6Lqy
8z+sbsawpAr0PzY7ePwefmS0paJLUYeFkFM7Fyx7yNFCkG7RQLhzpZjqa1PpK8rf
8LzBAQqUBHOMScvblUpClvCnM18Fw4xFFsXFOnRED22UOucUGeCim/MW08PWlcMj
U5th/0iQ6hDCKzBYOHOqDDh04eq7aAtgnFHUkUtk7f/8dVGy9xvMHncZhNrUVILm
weVObJSB0qwuCNIOj4Z6CUX7FzKMfGLxZVM3GuzCRmGfeizOwoPaR/w9NEvtrHMs
Sf1dc3Wi1npcBnpvsABqpF5GAA3rqWt1b2shw6FvIKoC3inVjxylQ85f+VbdzpRq
GIslwc8dswkpOflec3/vaveN3VFGKk8I4T+FIll1mYBF4iGXKOJsI/RT6K5EAczP
40n8uu+CXYedJWVnHasCmU9hwnlwzCQ57SrCi1PKGoM9hmjvsF92UC+CmhkwabOw
cnZvs395ibb/kORynAsw9/wODX8jf2Xvsb8v+xK3ZOOEWNpKOEPYUkgHI0US/IEt
cL+GYDu6Q724ySV19tJ1L5bjuYrAFghCKyVCFq0FLAOHw3biB/hTvovf48I9sGGh
DUeYXzS2QXVvASwitInZHRVWmksrWMQp1dY3mmY3AnXF/sakYAy9vTlMEfK1FCvh
auo8HgWFvwyUOVcXNE9cNCJfXDbO+OdvUF6myXvv38DKk4+aA3L9erN2WWZUQHMK
TNPySPd6OPAa8fMPVDzGHT1EPSnqSTGLuceohy2BOEEXVBoWo/MWQ5ilRt7JihJx
7y/0AE5ahLapxmEJN1IurpI+hvOmpHAiMJWNaFb6yw1gJODxjIkRHXFYRNTv2b+Y
UXLXexv+ssAwzv/v7RPI8ijA06fjT0O9nmLU6AORuMcxXm807PdB1Ns0LnomzTIC
b+SJSjQRh9/s5te46BXWZOk1712k9aKIsh8zGXhBmSwfAkQXFt6K26HMAD92hYqX
qi+LZg+cwiYTIr55vynpxY0HUbWAAchs9d5Kcp9GdxHzQD8Vf42oR1+NG9k8uqig
QIZMCtlJnjKgwVuoxZOzZL2QC+eXWSbnVMvG+OEN/iyT4IhHC7iSUoxfGQkL5SX0
wGmNnLV07iZpxOxnQ979v1Iv4aX7OnfbzwmMyIvs7oKOdXwbHrE+uGbD51ka1gn0
lgx498Jg0iuKrOx8/cRkM3gisN+araFnAABZo/6AxUi80udXwkf7cKa5jBnGwlSp
dFpXFWFzn2SmLry3q0t3PPdSv4i4dKKMB7MxQjFxfmY/bUbSr6UxcWsommgsm+p6
4z4jKijLlq7eQQmX22pPtMGEktsZhXYMH8XxSv1y/lmTtx8b4643Qc2heG6wBcTL
RC3nEMrZaDG+sLA2YSXR3x2xHWcGyqU8Vula6vVarqoaNmN20FvINHcDeKTjZJwQ
4G19IzT0G4VqQXwBWHRV/Zvrdcq2xl62TpvCHXyVJo4I9V7lBNZ4Wha481igJ0OM
WoEi6eSn8vuQ1mYY883PfSE+M+UtWWqjB2S9AiHvgTgHmzKMLdcWP3vGgvg/lyqG
JTnjcW4RQx1xsj7Az2FMcd1v5evcxZJRkND7lYbCfmlDt7k9qvu7iY1//GV+1aLw
ftWkXnBdejzix/+w234P4U9IEMpLGnSGOF64z5OrKLQPy+BmjN9VHgifmb2kjQFP
zJnol9UYqQtU3QH1EetkK8AX6enAltzsqC/+5vA2y1+DKYk7gqWjga+WuBp4As+b
32r2B4ecr1eXz6UcpZVqeE1QI6UED0lAz1XjNgdhKn6J0aBlT8JrBLxqnb2VZn/W
+DeY6d4nbMGORK5mCHzS7Ha+1P0apsvIEwZ+llgTyG+Bf8T0cOvyTJ1y6R24OUsU
qxUX/xuwzCUg359MB+mQcbhu6JHOwa4/l5MAOXudhz1BtZftD4B5KAa3Qj3Q1Py4
MkKwPXwWW2kibTxFbeE8JHnsZWxudeg/54Z/aofqXlQC/X7Bc9CRuzo7NlSLIspv
w04z5a+u5XqXPBEEtlt7q/iucMXR+MP+szu0NazooLAZ1IJnN74A7xctxslQVMvN
WGmGEF6GaAE7mOiIGKTJaTq1h/ON7Eu7TcDdkJi9pJ3VZqaOHdfYN1Mx4QfM/l69
F8MekW8p7mgjPhnsHA9liHNJnWbwZLUimsq0lQsNc+7jTTa3j84iAfQoFaX/7dZr
VMyQQN7HgAIi8AYOOnr/0369riSJfhgyaojJSqpYPcTHEyrALzQJj+ikIvVXsgZw
tc2GQc4gH/S71xGMgx7SqfQGypvFXOgexW3WeyJnHpClczsdOTmwb1VTR3pf9y58
912njyxskId1Q0quY9oqDofztX/BJQhGfJnZYykjoqSpj9f3RccdyeRsy0NGL3BE
A6CoWWkvASwD8Z1YPkahUxHyg2QF8E/vUtSAsZGCkOEc5pzC3IBFb56oGNcr4mdB
gzQoHSxWjVi+7Jyk4YGGz2vPIlmQZIHROGkzY83P6Ri7/kDOlmpm3Ayz8wWApv+e
oBF4RwOqkZKPYLqeLI0fbKTNQPee0+dlFy8XAq/Y2Ct5YVARycSt6hJp1p1zR6ld
0BYN9sl8hzQ3u7Hxnwqgoiks/th/M8Ufpm0rUppbOEG894gNcbaj5AM2iVkNG98w
FEBFv9z1SFlx9KoEJgo0DMt9WiuGtRlSyduWs+fTdWW6vKjNknUjjw6H6v8eJNyI
YAyEvrE1+ttrLfJJnSc2892FvI2tiA+RSo+c+AVQ4N0r9UXwBhfutnl+xR9RJZUn
+obJHX8EoVOEhY26KojfoPK3VfINzdXhbHJ5/ablcMEFV8iCA+/3LlPAfPNbai8x
uDt5bGX6WXsF7vxxr8xBhIW9HNqaT8OCeT5xnhWVC9D4PjLJohJ7bCSUf2VkbVRw
I7OV1lzAWSd37gXOGW4EthXvv9Fp1MZHTHqGwqjSl2BDtKOOzUxI8RJrJtOVVUOI
H5mmDUnXFJJY1DT8akxMh9CDhjCsE+tKCVI0QKeqcuge3/7jVq4j0WTqW6jnrNz3
boELdcEXPt9fAIUZFSn7C1G2QWn7Tq8AZu0E5c0v1+ZROD3GADQzLEoPOyku571F
Xe0G7WWDhKAW6GDkAu11YwDK7LWwKm8FEjQne8BqXOwVEVp0Ye3YfzKPoYNZ3uOd
bM4Z9BZCiHA3S7bsf0Khna53c7RjSePNYZJPVh83riOPB4MXB2d6FftC8SL4L7Kw
04PYdSPTxBbTnwlWJYEBuUK5lKGtjF2k7L/ES3nZEP2fXQiwogJtFo+tGJ/ZCRrh
hIfRsjDBMqEtReHwOO8nmV5u7F8ZAOvCor/GNEyMDP+7y1gmrMtOspxJ7GbE66AE
a7nP/ytsCsk4SGBuJdHdfV7RFDQ5xXEhRAiEsuYgZoD4kK/zPmzLGtzmy7RIV1mI
r6tIpCUgplhT4DYh98rS8m+T2ZLRhysm/aW4iNWS4P+qudX8BK9SHO+AuKsfwPXM
Dr18ge+3en+imBEaWtFeld2MH+/zCs9Q5/VoMRacspDlpvyQ4gS1xSsYS22UAy1X
SmG0H5G37Hg2R0d9uMt5lEV8vZW4bwh/5q+NoH2PBZhr7aNWwNQ40x6y8oOAFjqH
2jDf5rftBTDK9s9jkx1OuSz8JbG4UPsBrpN0LeUBzT4lHOpmkaUqLHv2AQcSwJC5
qP9emKidXysFHrtCoWj+/N9USs4PvmfNPIA1AfAnLWIGAIZOP93tl7o0UlAqxtm0
bWed+cnjrpL8teyltSMx8c3R+sF+tF85bfJnnDTFLmvxOkVSL4bPjsMndIEzJps1
YVfp8Wg1CJqwnhF/M40JjPZnuU3D4V4g9LnIKbpC1b71sdoOx/ZHNMMyh0VGePfh
vPRNgxBVJXoF744OyJZxyMhKGrvb6KFIVyPnzaWW6qoIwUmFkV3l+YDTT1nHUE0U
IQOkBD1NAzfFftdT3P7IKoIaQhjJcbtx6VJ++0i42xgWGGkOw6jXe6u7SRmwTKnR
xxEhSSJOYw77JkGCzoDpHgEN9eCl6WTAkBR+mG/tlcgXV9vMJr3Iao6sZpPtSas9
K2yTUW+h/Yshw+jI3AAQYsZ1gsSROeCCB8fQXmCYNiTM7jB6qS1JGG5eQq1v3ICn
Lhz+HcAQuiZ3T60L/cpeEvmoRP3U04RRp0gLr6lHptap+lS237YofaeQeD6Dkm29
K4F0n5Qf50TSgtBzEoAxoy9auHK/VwkJE6mvgvxS6HL/gaNbA+GKcNkshvVyJM/3
CGv02m2nB9GtxZ092OM0xMWJdVbHetLFU2IDQzkzZj8BBkV1p7N/ZBHvge3KukjH
R6NqDtrOXzUUu+lTdqFvufL+fYpQUNdc/rQwzHNxebrrOdnpdzlBXULjNIaYFFJB
TtISeL536BAmDZhbAlIwbMS3WikGpBfftOdqQkE5m1qsOzel5+EwClwNaiBz0BEf
hv1LfO6GFyIuAQGBtkVSMyh2ZDeKiFJXEnG4HRnyR3dfsm9YNk36DbqcEctoZIW5
G+Si0NrJnDX/GCLL+HT4vna/ZeRUcUGM9S/25tS+sRN4kIlfHjIGXKdG5RAlYnzY
fXO4pdGVsosk1JUYl2R4W9ihD3acQ402ZFyQSol/K3Dpi1yr5VOFvZwcVAU2tYzT
j6UoLqsftfM2Mbr6n11KFq1am/8FbkP6W7XOvd37D30EB/+WME17NpbluDYSRgjs
vZdSteDazxzSUnOiA7cMsrjZsr1uX1SGYhjYYSZeXCdWvPoFnjz3fH66UGUgJ6pM
sy/lZkgKWgAbkvc2umcNvq3U7pDO0F4doovYMgYV/Y+Slbyx+w7e5nMi1AZbIpQs
EAUuKay4nqbq3LUcqyUXpsVHxS5tzi1RlduV70ikkYtmDeI0FSdCyn2sRqOCXw3b
QfISoPNFIDNUM0TIhRL0Y5wTVD5Ep8cYG7eCTxMSbD7rzau8wxaYfI+SzEau/pDR
kBlWA+bXxpLgQJP1zpa0NSZJTBrCAyIgF2FjPU6oBS00OqpzK2f8jCbNKIwaJ9Yz
I1yO1qqKLrFOwoLTSe+doHxUjbxy69DfNMGxuqTF2l4z1n9LITU8irWsyTvHT384
n76aw9gnCn25rIay7L+tb4wHTn7Smj0wd1FyCWMDehlnknUmOJzw4gU9W2sUumx7
OBTehI1ypvfrqfcgkMlC9PYuMXofXXrSd9AYUrFT+EFEZCAX37kkSIiw3QIPFTpT
RP9A1ZQJleHbz5xF+A+Q8wAw/Cvhfso7/I7K0kXhZkUmWG7rgg6jEsL1dbW1561r
egRpZmomEq1S7UGCUIOkfvtaZ4wuSUK4AYdBBPRK78cwgCdGUuVukLqdoTVhSV2b
+3W01Nb0wo6lkVui6xaDFK6qyyVxVQGO0J/uSoo3974aphuQrtIdF/khLpV/Va33
bnjixyDarJm3vhyhkfyTRsAL52Z0ptwWGfXLuKNhPpARqz07adGG3Cveo5KD77xP
iCifizwHnLsDGNnYqN5Cmp87yLC/Pt0G/4xlEcCuTpK4xNA3FkcBWxBVrUz/QTEq
9jki7RQ3gwCBI6vJnZD9H0fGXfD3cFwFI9Hs7kZzsuUdKYw796C5MvIj/s7WYUv0
8M+dJTTY65/Paua2YOssjsAW8u0HXb7LVsCBi/3rlTFEo4ssJUTLOwkek6+wDyCK
o5p83OzsV6aDPzENAD1G4Xnoh3Q1TrrIxeD+/PJI0Cm4Sszqc75WGw6mkzOf4sM1
wPFh7tv9COS4dd2SUOSO85aGQixO4GhGBbFyy/+tyJdJlm49FFn/iLZJ9rMmsjqs
E1AO3qs5Do4IT5fLlNkNAr+VbN/Bg20fB2oMZ9RIf2e5xj1BllpyuxMOXYCEeDUc
k/ASxTcZIUwKF/DsrpXkWO+Gn7XAKmwh5h3liJ7HPDFX8nV0sQ+7xKfnELTHAeHI
kB0cmHZ2kucFgw3X5BTBw9ShK1ZH9OZLSMJWOQFhGu8b7XsL4NJuU0L/VniAam53
djUcS9AAgCbjwzilq0WbNSBa/7Xi0LOxedyNoWqEozZ++ReyjdOVJx+qWgcwVbiZ
emeiRPwWll3Nm9pRPTJGh1hE/ZY39wsN8i6gXTCX0NPdccVZdhiwgkgazDotCvA4
wG9Hdrq9XNukxeg3JS94LdLz0JbAwTByonDR9Jz0ny/HdRKIaEIylX6OQIlv/hST
9DmXXqyei7zSJuOmF7QCGxHVgwdKvHT3m+zLo3Eub/G4hEzH1DoBU8kKsOZ67YU9
yQWdhe7a/Q542eS9eijjmBkmye2fgELI6dw1fbWC3JVM0Xa0SYK7z3SEIASEFFXE
bZdSFhA0VgesEGUuU5/n8vVNKvmiUaWr/lc8bTkkji1j9nyRqCMuHTRJRpF73QSA
QXoazVjhlVnod9yfsV8sykBW2+RVWkXIwG3/LdG0iESWcm79K4vtsOY1wpSlGj/n
Q1/5rGEzy+yowdcwJ9R5diqqULuLuiWK6qulWrSlplFxe7R+Qo5zZ/AJlGdhtViQ
N0pSlqQgNomNyN4Z1qFhBLeND1yx2T+v/AwVu9JKp2+8EokZVgcnnfwcaFrzD6K3
6N6puz3/ZfpBmRQTVD554E3WPJUklF0t9zpyQoJK31briMQUwblrxEL1PM4iNJLJ
4WFoJb+UeVkLI7QyGCU07LidGjdZKqrIKGobFAk/WQwN/wXFsIHOU478YiJrDzZ6
zn+UlP/xjXwehcLImtT3O+OI8uyYSGxGT6phL1+KisbQzc14wVf6dsA2dOcTVgo9
5dxxqI7tT6XYKINAIWrt3TKxf1ZP0DcdQeeqdpqMJ9qSnlLRP3p96IqUsEepTw9n
lcKTNAuxL8Xj4CgMEmjIf75joGxGRy7eQvSqk8aFs3c8QYf7JpKh+sO1N3X2UKry
2VYSag84PgdR9zIyI3dMMS3RoJJQb9w7hmz3KoHBHuRR8PXArj2MlEX5tNILUDW2
he334YxK49ytM4vDXkZD+TXVH8q/OD1uwCMJrhMJbbTAUo7VnMgIBzD/51spYaVq
PfNlfVHkXnwqNoWuZcPx5lo3ocIJljmzmswBqnCS1YrbNhMbZLVO8T65GVji0+VF
BlnssR3b/hzMiuDNlH1Syvfo6rr58cA4GPAMb5d4vgt/qsUWOsH+UnMh6C7pgstr
IQKdjEy4J8kmRzW3NRCSrUen/HcFrZ+EjZXUfy4Qcg1WQRY39u2BmiP93Fi2RA1z
huAuwOyfybDkAmJrNc3hv6S2VMLNJZMF083cJ5WeHf6KLr+6xI2NKAirSj84YnFy
U+fS+umfRsphKSOmWbMpW4KsG+tOcLh3Jev9oVwMWxOcAYlbVTvsahNTIF2LYZ9v
lH93gE8MqYbZ1mLgN1hgs18j388uAOCXHS/3CsBQJyV004D9Da5TYILQjr1vBIvo
CyaDfmjkKlC5904fu5jY+whD+h3MP9tF+qt2pFNzA5Blm2XyMrZCAXd+osTTkdfc
vrzo4IeqJXE7tOPepTOJaVqfkBEtWg5yQUrmO0CTBnxPWKkJyjzflYyneJdD1eho
05nCl+rRmxzR/iJEco/2/U/tVyozrhpoaWNlbIdmTA+FpimedQVGiWcXTzoP3psu
//WxE5tS8MKUKTUhuq0BHHUP2L12CdjH04BNhkwVm1hzpcqcd17OQ6iLLkxIEcUi
TLgKHCyiBgWS9PLTiLEd3oWp/Wc9wsZNw5zfEPtFqahLauKBB2Cxwpttps0v+MUx
0wDYZi4dN6/wrFY/aR4qgFi8xbRuhq4+vrW8wZeQF7gW5UKCFS4/gcEZ2oQG6upm
6ySax0DgkKL5bdrs4Ywv3Ei/iUfj56hRdS1/nchBlLROxaNtopPwR7XzQYXBodXQ
E8xOUJonXiu87RKvQuu1IeXdeCyNeLlsacnI5X9j48W3kt5QzWB9JcstPBVOngL7
dgxMDOrQbiDt8PNngRbRygDMIofzTMzwfoIPdpZwnxQXy9/jbP9a+yj1WgIH9G1b
WqlpMNfvyMLBKvYnR/bxCzsHJWY+JlwWUe8U0CT7OKjRQwqx3RpWKKMfKFfxX9C9
PW/9JdAfGXWNk7toIal2v2/305U3T2lw6Uoe6uVPgdgoQCL4RQlfzqAXxFEE1Z+B
2t3lF21t5sW4oVTVdmv/IxjUPCFtVjgGg4Ko23NYfcvPZx+A+9HnXXYJ9l+z5AUI
bcmYU/Gh6g5hH30YlrQZ90N9xF5Z3CnWr+X2Bvg+X861dlDgFbz0TFP2x9Nkti84
hwK3tkbgRQ/4d+mofcHPfK1wPMJcAndV4AERxwa+lduQfZDF0h28w/xxCNCqoiDp
53ZobcVfRD4Q4Aok6MYZ8wGbs9SbbgQiV9QPu3DtYI2A1xB1WhiV2Y4aoBzmnqt8
S4ElSpBj8hCb4OsklDG7lL1BdeXCgnzH8SRemlmMNl/3oUJaqw2PgJA+NFWZFSQp
QG3eTFOtzYcH0YUmkqSRNpEHTOG31l99h3m3fIkyYrkAJ1DNkTMCjAbkZpzDfz0s
KocZqmbTlhHr/9AFFstadSFb88Ok8srnxAEZN7I2a8jZJrjGI/YyoVGJZkTh2Rqd
j4htDCVbLZV9jz/KSM5BCMcPIlNdvSx5IQEqjPwTeHJhxMgV6WKbJGc0KrKEpBYg
GM0AexBBFVTt3z2E6cCCBJoqbBUjUI316sLqw4VRmB07yOfuU4Rg9IOe7Zed8HIY
gXUaGptuS1BQjlc1KvwZp5f93eQdDUHir1roEUXSck14tq3UKMVTNdOoDMS8uJxp
63GdgP5cs9HCR6l6FDhymIBQefc0VJP7WnWuN2VsnvBZ5NP9ooRE3aopPnphKsQS
3LQuoowNT/Sig9o8sU7XDfzwcdZBMGVcDZ0rdVKR8Mhc7E3zBnNyCV/4r01g/+zV
RulzNJAYId/h2jl+QGVIgn5mzjtVQW0bJ36/yVg+jrVnvLDBOyeuRtmdpM9LC1LV
FsQHwFUckOX22sLfbYY9ISIIkHOI+b+3uDwQyDjeauuh7toBjy77VRNM5SO2InI5
e0X4gZ+QYFL7l5/HK8xuL66Qy4wmI+cIH9VprMqWbApraq0ssOXlEb1WNOvtyhtb
W5IIPUSmdUAQjj4BmpiVwTQUSUZcuu1heKSiHxspQGUQCFST6OT863aSflVC97sh
nk2vNLhQ3qCFIkK4zieiPhrHszMQ4vp8+KSnKJsYM7P6/tD8xVAKdGRzsB4WvWbX
0TKX2VcoA8RGDJaqjJc6y6rW1waQy7IUlSN6QmbT0mc9twmn1MGg9GUkO4EhJ0dj
JsxImDcFBpRZbAeBY95Ub8LBi196q3aUUfULgtLSjWE1SUjV6dpm7MUp2wanIu+V
l05za4865CAn5vXfuioeyW73CDNMPvtQIGqC6wJSPivmvPJgFqUMrmvSq0db7GJO
nT94j5LJnhoRPBEi0eqtyvsAqwIt4JPikda6qpcocegr0oN8erZd6CDAb9d0XLMl
y22eOO6+UPyD6Fne9SVy3QoK8O+zw6XCVR1gR5I6UVRsuHVg+D/2lXk7UjSlmrtS
Hi3YXmQbKuULw9YCFPMb8/WkNjyx3KNrtuXsppFRhM00IUyWgePwMnH0Nw9Vp/JM
Ekh4eu2kfP70TBH82RYxucu5DZT9RXWiXsam562nP9c5t2lZcUEG4XaWuXMeeUaA
THvB6m4K5g+aXr2WoqAx6jw9fv5Jk9GB5F5/xOZ5YvahgY73hgenX6teHjTJj4qY
tQ+vnxGUGZjhLaD95NbBVwGjeVA/bBHRNdaboWchn4LLg26yHnriZ7UB5GgojOzX
eYVCbaeerbofInzCY0FOkdNjlyC1Bd7H6Cc4SKkfSJi1DfIi8iVyVqI/ecW52BjU
9mDrVoXYgw2ivLRe/FLBWUHnJsYdBbfxbg+NJ0t0xdDTiuDc/ho3g0CsmUbjuLrf
n9Huo+2/pD1xQ4IDwathfPhHvX4W2zmLueukQZc6UvPs3tJpcbqfSVVrox0uKoHx
/+hrCoxw9e9G0u9Ip8lRy5fFFN4dQu5oFxl8bNHwzC+rWCBaO3GvbknZzyXHxAHy
TvtiZvLqWEOfJkljnygt/5NGfEPINqsJALP4+SsRZtOQTWBhCgGSGvxDP7O1UWbh
58VzI/fdZ8BfqGEAp/CNKdbfIz4hVQRFnidgGkJizFjO5zgQ7CWeUbCjsVmOzGpS
oTu7e9D5XUAwUGkF1YYVqVhisum2zt8XHjNODhxO/VjTAxPE5WkwFQEqs6WHndmN
KysrD20qEYFcH8qqnYQZYj/LkPRN697Fg/IXxHLAxJLwNcDSc4fn4F1m7xKEhX+B
yTdMsn/wBvcGMZxUeJocIv27sJKRgDDpKM9ZFCqlujw9MC9kXOwNkNsMCsHcx/di
XOjQmzCOeykrMm1X5mf1F2HH7b6uVbk11jZw7w9a1MSw+n3b/7ekKQuXkcryxFpH
N5fiHlFYOzLR+hCuXEZDY65VVlEfmUrnOulzQWOlpWzaaMEDVNNiyCtZWx5zA9hZ
OQ5MbhrFD7UuH0NUni+otF13cslIWs0qG2/N2tm+/RYXAWQ1s2+whFb6GnII657o
tEO9RmfzG8WP0ErrvVW/OznZZvR2ARajTDQxj4vcJ4cWi5g54IaFlK/hwrtJcYWd
lhWAx0a8FR/40olS/E0r9YhHePs8zoLfC0n5DHf0rDHWPiKrAlG8hiJqYj40c8qF
/UzImfQXW37+8P8OOJpB7zVhWZ0Nt1s8hJI3ngRDas6Xk8oFskFnimdCLnP5LyW9
HKQjqKiJp3eITyC4NPdMDvYvczIuEDgurVZSj7nxDkARS02bs4yOH/6lJfAHJaz1
RHINjEhedrtbTkQcqCkoIn+rm+cPOh6RqxDBiN/G5Fy4K98k4eDJ0zthWDLVh1Ze
01foBFKp5VhLrGzhR/yWpVmX4aw2ss0gs8EZOozVrVqf9ARRsXQLl1KzqWMZs1qf
N0037WVlY3BrICAf928RI8sRsL73Vlx6HJQJMVq+KTf8M/pTmoRflSOTlEcB9vDK
gr2dMHoZVAEOoofcIhy5Sebyls+AnBsgeXCQVbjy9SMci+oNtyyQVn679wg+gYKo
8Csi+6sXPMWt9fBW/MYuDHhWKucf7oAiwXFNjlMYzkXMk6vubk97FyEnjJQL1LuL
JdbFQjaDkV1hUA2Bobv64EQhcQB3/xbIgna0GciXhm3nBcfuO9ba/9LsDBwzMZgG
ouVIw/5giPEtMP6TaWof5t7qiKXBzWKUrQiYFxudG5yjBYk/2s6KoFaUTLas5PWA
MAcVbqCoUC5yedjAyyqbY4MuAsEvcZwa3l+I+/cogDhKbjvRCJPNfDjYQu3LG4Js
y4CA4Zlx3tJvdniFV6q3s7pyaJ66LmMTxjI6sQ6Q6ypM79QpoUZP4wjQP3XyUrXR
ERD8ZrKhttPdRDWQ145JleJamxFXdeP810gM9Rmd0F1TpPi0PP3OXVHsRd91mz3r
ADHzSpnL6f9qLZJbDuc6uXds3CT5sOsTvZIBXz5JfIthQg3PglGqU29VFtZ8e/Dt
DS0zfVC/jhTYkJSZ2EUzGn/qthwQeRbXtzngp6geEoO3Jvag6Sf8nflRu6gvzTCj
4H7L8Pp/Thu6QS492Yj9L/jxfj0BnIqN2uNCHsHYc2cYs45GpDGQek5dI+oTetOa
DtRNBVJEGXAbj9eZ0fJnJfINtA3CYeGyEqil5BEBQbzO3FWKIqcUgyhPKP+20oAk
p4BmfLAsOKQKluHz5N8G+roKykYRqBlg9gTbtDtTnyaRjsNBdvNPE5o5g1vX9dwB
iZNuCbhwXWfm2mlvGtO45LmKAg+iQgifVx0xQDUSoaWGDS8Tp+ObTwgJixkXNGp9
2GTeQB/LxugrDDn3+WZ1K7jaXsW1MzMUGHrS2SmeyeujeEtY1Y35n+u/j7+GPjsb
n5s0D4Yh6F4QeiOPwFV9KBPzr5AAl8dZDWR2LJQZQ0f1bmGo8bDwZ0tYC9QM8XlW
zBay0EuP6kd5KfS8P4MsoSQybWm1X4zpRW5wWzEWoNkNKDRpJGU/CshyHzSSbMPW
5MPS53WxjjUqsm0YPsFE3Q0EptGQr9Bg5rFTa+c7f0yuNFhXRAf3fiTOd/a2IJD7
PNMxpDnaGBjqPEbPI0cEek/xD8N/IynghGBt7j4ciZFqH99tROxeErL7QWTb1wyN
ywozV1U7a7A+kx9W1UUUnLWVT0/qEJUIcbwBHni/HWeRsx8I09ZQwYMT0dUy1vRd
ENLKCui3uahqU/EMVZeWJHJTaPMxNY4pf9o6pI0qiR98lVNsDKoyJjZdzkV9zu+F
tRJ7BZrMq4uEVVqCwZO+DzX5xnc6fkJ4ByTuvMFlCQ+D0mAW+qdFH1JcfOTVT5z8
LMrvhiJA9xkQj0BRYK0Jm64IHY9Ja9/KQ8KW4oWKx0ihkvlHDp+n+lDaEf3/vGOH
x/JVNqEbWed22whJcoQLVqPLtabuWOUC0Tnlkwg4Bj7rv45P0YBn60tbbVIKNyp7
+ucRdISYmqyi1SmOIhaXB8zcZTTIQAAr+8l43UcJOaY6vY13GKy/27JVbwDW/1xj
3dqNTJUvo+WTrDug9r1x/WebCH0aMrcqbxw4tHpEPowbExuv+Und0akn7NdkBfO0
YZfdabq0j/BtiM2TdJUSmCJY3hjchcbiv0kXdLM8CjSg6dwI+vxNQIDv0LH0koXK
mutNLwK6BnvDOTWC0TPi5cIxQx0IWVKlGoDVvRwu7TBBFkKQRxLROLyMXSYWSvUq
fokNI5gNbIeIFHHPGQuaN+AARaERI78yOKwE8oUuKYLCr7Scu4Rfm6hLTdM174tK
PMjpHAOR4zCtsPsOQ5s3IG2HUq2LBjFrIY+K7ylxS4FLXtkFzvhRwUEhmRi0AzJO
qvnI5RMrZgc4odSIol/Nx9zCP5ujJng4HiP1Ppgl+9lxXXNCQF3p8AVLuHHnlOtZ
CPL1ppMzLjqvFc95uL40cvOE5dCS2xspC/tw20I+1q0CjBLxtG+G2XYuuh2yrmO/
nOWjT7Iz6fffYOerD31sFhhcBGmNrXQNBxQT29s9WL1j6Zg6s9tBnLl1ZPgxgYcJ
gYbmjwQ85FczTt+Qq8NVTKQO4w+vKGVrctRCB2Q0fyQqDkZE79OIefglDmnv+IaH
tgJ+6URYrLiLWL720ecuktk3Voc+aBLG4zGVEmifIGmhE3OwCrEBhPh+e/vBZjRc
w1GFXvurj+T+KyCuQD2voMKsoKq2EGCErWT+wJjxXAnOtSXEgVCf8DaK5RHljq1d
XHyhgam2jV/rX+yjpBMzQvpDGFjLihv4btf3BSSCnxzHYK9HSl1AGhwjqA60sttE
u03JGxpPqVOpTyrvJtmjC44lDtjY3NVL5I5XnBi1TiS2YsfI/cAHbcgx0w5EPyEH
P81XLAlSj3+v9IYIY5lkNzMmDysf8cP6rtKuh9Ne2G2OcjR9AtqBJokIOk8Ika0g
CrjTeUgBXpjPHcDsiZfUOBt3im1V0ahx+MZpKTZv+8fxThPg8enDzGSEAZDrtnUM
xfWJ6gnCprxPSgzdc9VlDwwSkxHlkFZy75e415HoISM+Kq1lHSpe2i2y1NUaKcvt
rPdo/ZRzXmO/0JXquGD/32oa4i5wi2WNT5v2vu5H9vCTovvAuxPiBZCA5ICD1Arv
TP+1F5entILkzoepa/46D9CBw+dXdhxRpJZHmdW2VN6UaRz8fF2c4m4Tofo5KQ6c
+2T9q2HUUdLban/hB9/ckUsUhGxNV4hJWWrudetepsXmHvtRGFv4rNzOFK3JTUr/
Aauhg7EfPr0oGN1gBo8W41eDSzI6ndx+0ZJx+Z4QawJRYo4lhebEHF+/ilfjp3W8
GqSu4mEJl8cu2Lt1irwNwprklyglLYeYvxkMBPsiTbw3JuAbbEizysX2Yq+RJ7nh
yfVD9N9dkRUxuFTVdRj9OEqzF+a+te7qza5eSAWuuayYvIbBAR21tCRO6NyUQsI+
zm+IVFsc7c7MF0KXtrxblyxK+nkK4Rz+06pH7g1+xNJ8SZb0/Lc1EEfavnyOAJSD
kNNdOxtdW3Xfmonx1UUaajkSRXsZ9NA7JAbXXUMSGj4mrXucTGEnXdZirMzq/t7S
Ujmb4VofIJ6pJLiOTPm8Od7KaJYTP9W3NKH7azQ4Efx9s/s+irpyurafkWgFuA5W
LvPz6azlvTmg7NRUiEkuxcRV5TEExKH+jOqAs0/TeEKB4dMo3qdjH9fniwtwi/yj
K8SNk/GSy/U6U9MAZSzTwvfqhzM0JqKSyRrUyigpmahpow6IdYO+Md8S60opbCyZ
FqSF8VUkPC/zWEcZGyNuvordJFsBdEP/4zxZuKCDXpd6phczeVaxEV4QGCpW7VyU
wZuZfW3ztRwHze+UFID9Ui7gYYummVtjSBqOYY10PTzjE0eDPTr0XS99cyYIn1cP
I2Z9L3wKyVYhRCEdPjFIfnEfN1arTTKuglLDZ0kkQmIfd/lcBBsRzLOXYc0ip1EG
5QsJt2jrDaPgWEtHcoJAHfyKmhsNRi8ct4N7Vdj8ypxrCgXJxQ6pONluzuEbjtFy
Y3AfqdJy7dA7TmFD5KSg0qhQ1oVd4wDOn2Pm7xyPRXlb040XDob8x82jm4vEvZGI
Lhox3gQ0uD2HzyQYQ7BhbyGVxSUmAchQysh8zaP/6CLa4bKfyC2aPiKgRQtPlXph
ci0nij3MrbZQQAMF6vvQlgiixNMzQliuhzm9PYSeMVIxOcJgWw2JlqjOC38qrmg7
6hBMxfIW25QZ7zQ5Z4AtJ7rU3i5SHkSSdBKSAxdGb1kTPxTtlwwfFH+phrWpO9BN
bi0Ck3mcnymdtwrUgZkjsAEONmkOxw7GywJ+Ku40y0zV20a/wsqrgHAea+EgNpM+
zCuAlBzlhHoWnk6tR5jKdq73JxJwu4uCzKaIyzzutjYUpnoLX+YvRxYw6RY1Us95
6xBRL6bDKo7cvtKxLH0N+EpqpY+4TVs3b8i3g4F1HqWymhNMs7lV/Ut7aZvO89GA
hXM1udQpBfu3uuv3EeOxSDErMwVd79t3orS1tqZOy+GWZcl4TqYT1SesiFD3GAwZ
TcvkUW9w50l7lPAbY+VKkiMWt5kienxKwL+pUL4JT39TiP5msoQ7RSVch0cf70aI
tRIJrridrsI3zDoKD4PtuxRPkJOv3e3959W2Nz6vRzdKZr+wNZRsgJfuIuA3suvm
wl628M6dS5aV/VDJZ0EXJPwtONz5bJmS/7RPlKaD/B4IJJeiyoojssxkdG8VyXZv
SCwNo8dJERqjRBUKSh9Xyd9vCD3Jxtt73DfLQtpppu3JRD5VyB6R1WC8ej/Usycc
rQvsSZCg4v4a2PRZlRK45VcWIslfP0c2ySRg//sXDXZvJlnPZCJgNADiedMLzJEY
MENtZa/tqMJeO8M+b/3j8sihIGiNjQTtvX0Bkw0y/13h2aNR25BmFSSYraV9vowC
L6PKLIByaP70o5i/404lJk6nkv6S5kSnx6+KYCVPWpVXs2YMy0maS4QBh2PFJB7P
Jv59Hk9WsXIc+uj/On21LVsoOnFbntsvYCcvn04qHkQIK09iVMgFvJQ2CZ1WCPRs
v/H5NH5aU0Mu0pnyRmIv/NxqvAHaBYMPHSI2sp9oXUWzA52xB4yKOaq21oo1g3Vi
k8WoNefCzF26iad2JYQ8PLLl1q6FdpidWNH/yPgRqr0wzlZ7JyxaqJjy+hElgauF
xG2XVueSXjZSg4PqapPTtaWU4CO3RA9iTjkJz2UiJRxqjZfTgakVSjNfdU+YReWY
9ERRB2oD1TKDMjHv114WdwrTbv0hh8v2hxCnV/JF5WRmSEZblRmXHsbIHcLouM7p
LEyoG8yN3mjFJWAfwaGSeoepu5w5swZX/UywYaSUnPhs7FtFkGASpQJhbZ2rBZY1
XhWxnEi4XP+Aw7lT2fyPv16BIsfqhDimmUokx4n4N/AqZSq5vlOueqSK1JApNAyg
TXCj8j5Meudr6yD3tsGE27lDTxN/uJM0kgp5dQGZyq8fr96HsGawQxEVlorbOok/
6/0sfnRZ8hJdY+gvw3fy+e8zk7dK0P8W8tyP3SCT6pt2ohYmNfXytUll8K5qX8MV
fP4iCiJ4J8pMa1+VwQVawY4Zmu0m6Ucymdh4vYv5XxqjEVv4Ep7rMg0g+Y7pdK+M
JP2DBXOfaVtN45xCl0dO2eSj7wrvY0tY0I3/mmRrU8Yh+SG7BbRDzO62EiLbpf8V
EMdj7e0hEX+RkQVbrQ8h2QXL2tQDiYt0CO+nso2HG4WHxa6xxbDzoDMoDlyv0NQ1
meDKgPXLRNVNY0++YrFlINEhKbxJJIsPMyNAUxTb55uHkfze/fanSMszqERKeivH
kQCTlf299kWUzT5NskIjhaR22lH6IdE71SMjCGKtu1N4D2nie9LgI2+75Mf64HkB
QdqnGyDIsHxM89Nw9obmY+4N6vzJBuqu2pIdQpM3/iUj6POG/jKhUWQ0N53TvR7M
yMxjlc7/fwG3LWd2prEjKgDBomdtF2QkVN+uokSFxlJUmJRQEa7v+0hodgH5L6fj
XsuV0EH00BSFb+asmyz2VXtIlR4k5hSN8jluoKhzh+Vp8sQ+RSuscVDEgflnK7Ts
Lregd7lZ9I4qifCveYJiJHiefdq2NWVyGk/PAPe4JhIMeuk292RoROt193SznXdK
8CEwO4pLNaxmKiB03rcd3QzkA5HiPbsyyP/bSCGLUH4xEziT5xhdnDnBnYLWCPqT
SXBlbuxRaFTgaNCPImiMkhg6agW62/0NnRxdvwKT8V1PuNvIzPyVgVwnuxeiz9md
hxp8EKe8J0jjSTEHnlMHpkYGW3N6PkmoYHF4Ql7+xSdEAbVDM9lQskkzEIg2L0vs
g2KXiplz4KvFnkl+/eeTB9QS0DGA7S2OVQztH8tWU1i94XKcH5cTyVIXsG4nwN6A
/LekUsEar5brnJ9lM4uWxmPSROKXdC0crsxjlFJ5HTjHDelA3+4UQiSKuaxySnQL
Ldi1p3sE5eYxROyv+KOSCifk4sx2NR2XM/doY/yv7GOTtiVW4KrvKfgZ35Y4j/DT
KRyi7unbVC/tEWGYM+NupFpXUao+jFWXLQb8pwpk4I19VUJvSqy/BuRGX1zyKJad
1ijPHLJtR2UvzJq8k7ZLmSom5Z3TuT5c67d2Gj6H777J+531qjFqYerBa474WM0c
URUBlVufKu89j6NfgcaqoigN8AZPKAvCJ71xX5bUt5MBV6Nv7a/Ltcaiu2wFc7Vy
E/cj23EeYs83YfscXkKyMyI1s/aVwTuz588zd9GNp3cX9ot1j3+2OKsKp9+Eim79
+5uJGwAbIL9jdF9J/jiy1RJfSKBwCMcUyh2SbFMySk9Co6vvAXDFSFhT+fze7gTx
aQhAvAu8vpgnUdHZuHjY3chrR4Q93S3k+YDKUNJVSKozHt+jllAv9RDDwLWWpWPl
F6/rbNJdERiJtw9ZhLA8ChcVP9jzjdumjVlQuy86mULo1EgjquwlvAYidMAnSpM7
nSr/Fw/AIk9o0l9HI3yPA1Fa6j1V2RlffD9WtchXuc+jM42sO1Pft5nga5IZk5TX
IkT/xUYXXtnf90yf+KzOA7QS2EZqxIGMnNrDqrD+sveusQIqO65h6+9+mrtPy4/I
yKiF8ZXmL0yLcCiOaT4I2f++xt35qLohhoIp17TMSgVT6gNupxSPDR6Kccvy1FOq
0iCXuQx/2BQNvVcqN+VeaBktB0LkJRul0RTaRnUQrEDdNQ/rSjHPHpDR92Zh3xBP
dPhJfP6ri4HmhkCiR+5XVkN/VrjgOTHCHrQOMuhUDeRVp8gjX3SGaswHiG3gjhUl
s50wTZKvIc8HEvS/iVUVoT/lcHgqG6ucF+NpHYnayrQH+XEuN+yrvnfasrWxrJW5
YcnAtFYc8l4QFjKh8L0kmfj4SqUfe9RrpTeMWGVbgyXGDmtgDJ/VCM+xb1iAat+C
SLOXGK63BVVhvYQtRnhWLkTJNbHowHDG6B4zVhKwOyCR4WsXej4ZI4jRL4Q7oIfs
O/aJQm5Mk8HI7DzhJMYTyWV+SkQ4aJJKxxM0o2r3THAEkCqN7+UFpWEIwoyuIzP7
Tx1i/XBMNj4C3sYd4mbk/7R/8ZPtWPGLA/j8X6d1/y4RpLhI5Qi1cD6lvwS0aBkt
qXKgtQCFdFbGWIOMncwzxXl6e5hr+pXw1az2UvOyDfJCpFwAYnr7j95iQzhnQBNU
uaBHFXvKjQ+7h01atCzGpfPdOpWRFT4OPgpL+2rlTboPaZoYcOoKMfPDaYjqL3DU
gMxxJXh+2DYCWRlobMosOEKTaRpEbqIS1krdV7gsm6PazfwjMtoO5ZhVeNls+KQV
3QedLrGMyF6CCyasXbDemzvjYYondjaOFh0U6AuHkpzm2eGMsJQUCPHTT7GKMWpG
xS2kbeLj6CLD17ictubJbFWOc4UaH9t3E/Zif9VjFN340QHDf7u1DQ9aZCZyvRSP
so2KjZFfqg1DYvG84kHpBvsLcNfOQMD7reXLvekuOfjl2idAIqMB5/Lq/qq9zGjf
Kc+zSbZ/0g+wEgDqA6QXBnaW9QpKIRnQFfW1jsxQxf6CdaiE3RlG6jLiRNELdTxP
vbHpmXpqooEmajSRJx8+1jOZN2EPilrokofmZFnFKNARmP0MKc7HTzY9pv/r3I9Y
mB24qyPUd/mETsdQoJSerzAcLsJEAAfcLercgoTevEaeveY4ijLrpsp0pJj1PCHX
BBhaIuv6N8faLKx+y9WNvYA2QzVEUDvMhtYydmXMcMUf+FF5R+yQeHj+ZI1uBWQi
gsogNP/bOaF0GbBnomGG0NcsDAV42Z4UY8DtDYIsrWLVA9iVcgQMNfyDZoR2xmh8
xUeeeNhSuBeXaFGxOEGKgt69KSFAUjf8JpZUKh6wDjmOUf335BV9xxWRiCY6JflI
2aqRPORMTJ/gtcprKowkhVBFwH/+YXzvNx7orlIh04qmQbNjC3N6oWFXO/vWzxF1
kVoKS2a0/y8bpnDWXYUtjHzY6/c1ifedkZiH6um7P0X73aM4q4mDQcPWWIHYIvrw
vPOcJD3qnoc+3K4ui7gyvmKi6asXj6taz/lTrpSkRsOuEsoQZ43WSaDYMxoB1Y8z
jMYkru6vLmu6z8BTeXkvSZWhHJgjd6bO53LcWp+EAUm7Zg/hRekUoaKjmmHv9JWH
qt/Liy+BB4fZFmfCzeygpqyZYh8ERmVJsH7bp8Oi4JSf4s9D/JeWKm2aPFFhLW1k
dVPOMSCBImGwnlmEEMx8i9thJZQxs2lMXdsRVqU+AHhWyxQqXSL2CScV+ReBLpVk
qWxOumWLON60kUQhqngxCnSKT1B+7T5TYBCjF9Uu5KDeYsaGbnkvDyGW5CTtM5K0
lquVK7fgtti9nwmfgztOz0ZTwW1BCuy+WnQUAU8OHp/t77aGdZ2TgjZ7Wy1KhCAm
u1aDQkh3Te5gLTs1zWdmAi60IOTO/elUgK32vSu9deM4t6P+/8fTbTxlFewWz9hY
YGCwhmCzxLDbxweEiEl/Ojp/1SM2acg/FanX3M5MCvnkOdaHILFVw91WhRSGnbcr
H44lY6wxO92e+6lHhiJ+nwcTgHXUQ7XAF5vqTptthrU44spE7ux3pxUkbRoZII8J
t0dgjMg7IQ+IKwflCW1FG6T2VvyUZsvniGFSUFDDyIaRNJnxgE+8GtDQglHPocy3
fvsi3CZOG/85CK7gMynaRXVN81ObmZnRJvDaiRn1voMyN/SwdrizbjiaVZVFajZP
fulQTHJdL6iq4YQ0uYozaWEjHVF8k+bIFtspfYmBM9xiotIvv7EdJa3QeriRbReW
V98cIrMA1blExiY4xdRwh36xrp+jsJOLYkCKe6Uh8wjcXvz8qRnlq0pIVeh5n6b7
j338gTG5sU9oSLC3ko+CFxzs6jvvP+60IkQ+7BX3HFWX16tY0n5UncmT7bgw7sZ1
UJlRwRav1RK+zPJFD9qYb0nxbO7eB9EitbOXe/BuRbsw8ZnBWpBik0T2fIwpMJp8
afaK6oW4iBVWQ8lsXPT0GIQPMEfnhpikhgapqpNifnN7o/A7oeG4qI2OdXfzgh6i
HG6tlKqKvvc5BVMgjKCQkjFzE96FLK2CuyxFIVlcdm+tnadYvoMQl1EOCARhmZ7A
uXgtfgP6AcwJ6+TyVGW13zEDZciuc5vd7ynF71Z56Qxwg2TJH/jKXndQC9wVK/CQ
z/ckTgTOZSb33WchVoqPI4422hYMulUWNT80emUIaVmkSLDjKgluXbR4CEGGFQrf
s8mS7lCt54pqdcNbPSMqH9itToa0EvCIq4UKCEJatAmUJDyEFoJPQTY+6QIrkNIj
qYj+OTMNhnb2ihMSb/0+J7LO95PzpaiEORc0KPgY2WawOwPohILaIuSgd6N/lefp
/KVqn0xPTXf8YRiecGm2UDJAYoK7wpw6jH2PNoG5GF9PkofOfBZDIaP3TfisPnQd
W2Rm0RIL6CL4nvN+6NSzPtjFqzr9gkjaVK3qluRuUP4roFXW4u5uU0QvjwJ2Jq8A
XH9rJ04KWM7UMDqBQQH6PrM7FwdXFUlGZKUyH+ypSavWnfn8riIWyWA6tNzR5Wn8
uTX3rXaL6UxsmYnEAteGykKwx3HmIf5wvw1hdcTDFG8egRL6vlQNTOAFQ+x5haaA
ucDlGWGoDfhJ9KkqjDM0gs1U2OM1g/QQXGApnW0vFxxqXdyCDRX6iav9JDafQCBt
z750pO0XW+S0J2y6tNt/eT+3c0hkrfOSSz3j5sLQ0VDmPEuG3d/8PC8EXizl8O9I
Zss4G6UVt3UPdPiQVV3ELRSDwhd290GXufhiVmYwCnsJrwjdIhfPDqhuuKzKvqWo
ECA40xfcFxw08Sv1Rq9YZitEsXvLCjMHr4mlmvCWtqPp0LyAWA5U8uavdyK75mqP
+grR7XCy1YouN5ST8vZZKySxsR6VF2NbJcIzfDPMZ9349Ph2gLDSWztJawN2orhb
SyYWpsSEBoCqZrL3oCYMnzakJRQxdIvbqFtQz2xyKgRaSc74N9qHXGuFx3Q4yytc
ius54EEZQuC3OwQZ1QM61/k+24fC3FH/0WskDAN+2WQdsiRKR4soj/rJM8ReLaQl
j1yeFKj8adVwwOQalhLh/0HJnQ5tqCOYqGEdEV64dzBEw6K7SJiFIABnrrBzb/5c
YEXLEqvkthbm9aFbZaK/gZRxAa7D2fV4xojMs8LsPuKKdEpv5qWmCvKKdiTOqtgt
G1ervH1DX7dsNm4C1h1MQOdw71e25YKyISv9ZbmjFauCruqYsWG7InortgNgC8lB
CnqY7RWsfv5MRGeNBu0NrOvv74YVDKDYNi0f2CkxaPtwGuFB5qseOQm6xKJc7XWz
4S+w7y5Wd/OzXbTqPFNjizN3XrZo5l/usfceX7MoK2cjP+21bLxz/7OCWKlk5nMH
7XpXAslj91199Cz1M106CQB3JZ7uiXbE9klw43+6R666XfqiNbrn4FL5EsxxOEps
YK5WhFJyYyZiGM46G3nbzjO4xFDeB/gbXHmN4Qx37baB4k7Efw3RYvGZ8OA8muZ9
7bY7mbnRf2rJ+9ux1NQOAKRIWwPjPvllhBc3vpEHSPfNsjnlWaiiQCzjHZWE+C05
RL9eqI8vH+Z8wGX2w4l4DRytpU/caPhNSilwiDmvboJGCzQIqqw1kilHrfeNm1Bj
UUy0f8sOdTe6kjwvb/MORsMzLR51Ftjl+qnvWxr8VOzjJq0qoQDqHctrEDQwJ3Af
g+AJDblqH+jXu+mDAD8bAwD2ybzZmqNQERiFae5DwUDaIj2tu1I1K8hAVMPr8OeB
hDIKx18aIVCs8l8rP5B3G7InaBduuk3Fn51VM02nErsBMRiAe0DwzflhC31J5iQj
hYLIW/h7DNAjHj9lykq7AQ+vZicue71Qu1/ZZtJ4tKzYbR1EjGjt138QOb32F9Dv
h4m71c6XsmMBYuzAXB7b/UdnMTq8N4UtbCA9yY60QxFYgbFNPZ/FncX2D1EkdvY/
YhPhKzxQUY0k70e78mX0TeZm3VVETI5Q/axG3BKt/6EhPObYU9WIL6p2jBRalJ7h
McCwn2xIuvAJY2zRuoY0oWoIYuCWVC42gaRU56iHiBdYHwKJZhwLsuN+BPOxCCUf
sq4OxhhMRxYCi5yv0bjqaCL5X6WwS1H21WKf5Z+vZU0Z+TdI6lnAA749dVs1QI6t
p35Jz2A1qN57IrruQ01GEGSSJVHZpTyn4n0ac/RH2812ZvyCjJ9EywShf4pbVgL8
TJzi/341aH2P7ZIH5j7YMBcs6keRiXC1flEs6M4Ro2zk/7f5mnOGFlQ5bYtAICuz
IL8xxTvasjZ3F3m9eYJjpidCCSoAtEddC0TBKTZiwOqxhTre5cBR6Rol9xTfHtly
6eOVQYS+ET3JaJ+lU8u5GdQfZQYJcwLmV6HqyAzO5K/dJm1rHXhFxYGg5tthzIgJ
2fWSHLD6XApJv+VY2kIzjcy76NWFstLMn2/+PCH6dsSjucCrw3hiJFItbNE/PlJe
4ZskRne3cGBIhivGo8QHO+9OTqmypZd3UN/EOU/NOjhsZN9aEwUBUysiYWrKllBO
KlgOJe3aZrMpy+GzyRq9uBE1jDTO4Npg27V3pbDQk91yQf2MYUa7O94700vgcU3a
+quUxwBlo6FSHCbfCAwUuTvhumtHgGh+3ANbUXj+WIC7mTgTlfWOH0Fo1kHYhSDr
TBAO4DsSB/hsimOQUn7tDK+aL/5lAR79LlwlQiBkw/P3ocAKb0sV9hphkLHYpZ/w
Eh03lqiVxT8hMVEymwW/V93zJ2Xbcmk+TDVWQtzg9PWGQdjCh1mz7uhQ5ufb/SHz
T6Feya9xQQJ0+s+FkAGotBzKpUWlpgOu6ZAblsVqFhJcCenG4u/UbZPcn9/+B1G7
zkx7WJl61GuCH1n4nEtnvjYpkh8Y3wqVUqzhFuQhU7aDJSMPLLTyxY+gZcymtc/S
AywFyXy+xGyf3mUe4XMW3OwQxY9bu4E+M7moPKVMDz5j5eZEBWJMpKBetKT+a2da
Ta5gUy1EspTIEMM75ttfoOjiiIbmbbhZVXpG7YUnW6CiAQw9WxBU4xVVGXPiEub9
CF1Q1K2UZL0YPrWneXYXLefVkTpCR/i8G8oYbhOg5B1bojdQwpBgcRTYVNDIYkCn
hjYCxDV5Fx7nT+vcCXv8d1AN4MLfp+yG/7Yz1GMfBNGoDbjPb4cNjLvpvuPSXM9A
nlZYyof9bSK1Ti2te6mmDwMGRcHj37o+SLSDmMHRMGQGoqEy6RnU8Y7a2OOhETiH
5wXImtNnw2gJXVpA4Elb0GbX7jRnyRrVnito4LdBHaMYvjGLa/o6z2ZIwMrCFgiO
F5DEKwH7Jlx68tW2II7LvApeLXwg8yPucWeAgpGh1JPrc6+6So0+N8j+ij/PYDQ5
LsvAddoPwPqpHyUQxxvMBwVd21nvGOr60Gc00mOwbhxDVKTZGGT8eSX9O4cE3MSQ
ueFZuzibbdsujEoPiXNGXhN0HRWU5Wp11C0NcUYKlcFM6mi7MYTahvIHpimp7WXc
OeqpFvMzbh57xuxYduXY0XRcro0kWWZ8/CTkdsWySSAiE54xDKfNQEUPs7jyPCjz
7Fk3HI5qnhcRvy2p6aU4UPlQvUb1F7Q9MxjQJ2TOrmz7g2j84mn6UAZMHn7vsZWh
aCw4QS6+WPiDMrxmaR/rsy9DDxMRT4AAkm6CKUTi12U51wwIcPzoP1u1LUe5RXlr
cLkU33mqDup9rgf3EbHJqnlwaEXW0cv3sT3Xx9MSF5H7QjIlBHrlNoWd5rDJeqOc
LXSZhM+S9Sh/65IONn7or24jmh9YnqUzjhBKJgjdRtwbqMZ1Zsyz0iEtUiJSyYAx
eqTswu51KEFUG2XIhBhEy8xc1ciaJEA0TnGtVchHL6KSnD9KwPQOQq/2uHqd/bZJ
wTThWftKdbhUKZBQarXC/fNgvNkVWVwSYji8fk//yR4rrQPSDy/Tw01HpAdjpM0o
0er2zUcQe/2m9lkZbrJ6VMYNAoQjyWF6q9m58KnGpmZYjxhfHvfb+CET4jlq8rfr
+KDF3BVYtrg1WY2TXQH/WWEkVxyGwX6a1z3nBfGPLNF9aT9OB97UCZ54sTpoZe8r
YGwojtLOtRgaRGGkWzo/yCTc2zmhqe7VDvTNoU/+V+cgXLIhSNAtfJeyQVpyN27U
sHTA2F28mhZWUMwJ5FIi/XgQkqiyyrM5AOIUteEYTEtI6V55aZgfOSa74jxfYjWT
nwdd45k2uDK3dhAUhuGwAPhylSAtfoEFZ4gbJGUgJsQYEDfxg6elaTqNJKFFAUnD
2Ud499j2beqkvXOuZuEZa1rr5yoK92EAxpIPuGCnlqAh+UfShvp1TKmvDFilC1pf
3RZeZnEIkJep+uUDSpP+Lzs8fuw7eUdW4OtUOo/gJrD3p364PqMQhA+1wAtpY6JC
AC5pz9NEaJaq6zZuOXDHocH7f9KD4j6VvGch3rjGsaO5ayEkJiEfzRLNE2FoIDWQ
tQBkV8IGl01KW/jgwlewD2o0wOB+Yq9BKwaw5v4Yys9j//ZInWjcGf9dAXjAnysF
hW3N8kYT944o0AS1HECn/l18Q14FBOWQs72iAVhoInvO1K/5hR1oksZ4eiYQX7ke
oP5WjBCzGwPCyqTQq32H3lTKcDmj9hDNgfTUjKAWSKD+sA0RvKnVHhFkGz7kzB2M
F6XArn+xHv+kTrVfWJRuRMQWUp43ApDFdEZJ/zZDFnQlz4Zzknqs7jKaSD1SkTsW
NzNHZFzNBwYI/q6SsDVFTftib9OX7Hf1Z6yJQc+HYQSDkkPWJp2IC8IAkk9qV6T5
vvvq7TZnuxBQPwTlx+CQPKczqb9TiGVF1zHBPrrSqN22E85aF4YzboAeiLbqGqmO
rwx8WrhD29syazDFnZ+YJuN2PfSAh5W0YTe3wDSAK8YZlf4dle8PqV+Wdsm6U86M
TbxE5E1xzt0n5dJKqrwrM7hJlrwfITNEnjV9LaLEq2uKgxJIp48qnOy6JWL2aOcW
BovNXPfdIGBV+8MrtmKcrXYwYE06lqJLP33J1ZaxuytRWmFiDMacr6m/Kr7H5Ewh
a+GHM+npFtKTwY2IK5Ie1fwuY3G7RaIMTWx8C3/ua1c8k2NpM4F5tVmnz0gTYVwy
rrdOnDogi6tVuXA9JhUBZJSeVZEt2CAlTWbKM42AbeejaL8MLit86v3dxo3xtIHh
wRa5jXiCH7tutlgR85QfovY4dAclheUilpg/EC0MuteIO56r30E85mwCSivfRAhr
o2d/erC81Gi1RpR2IM5vZsWzEX8fMAZEKHt1uToCb3VKFYnLQG0eaFDmNhjm9VQS
csMcwydhH0MKlqf31epkySfGsalSuVQtEFo9YqjhWA0Gyj0cweFsFKSIXbZro4If
nJdLqMpdX/GNIGvfjOCVVhA7fCFDYPFAfXxrzkoeI6ez2S+9XcHvlW6w4zZ+tNOr
eXiZzt4paSvN2W9SAq70GXcZgf6aIC4YhxNyBk0ovNvuO5+tkDQdi0Q0fCtAi/jM
92tng/XSFRBvaG1XDkTpYPIRpUxzusPluwuPjOwZ1V993omv7uLVXUZsZqqTrVZb
cQVAWu2w8IIm7fwhjG/OilwsLuhq4nwIwsTyOvNkkaJqY2A6FTwTn00Yu0sg+COD
bq4NXSQATVk2SHcSIL5ZACgE1Qc0I1ruHGREyrFbsRZKzFVh78kkTv1WfHugeyEq
e6eng2HCqdFNwTBrBF/8AMjE0mqbIODms35aH58mYMsiExbe91U7rpbnBtwP4M8N
qW4dOeM+0lm25ZeVd/PftkYRJQ5wnJ14ICHPJ4oEBhEsrodoeJ+bfMI7CITGbkSl
QqVk7gVan/f49oWCStSPFTB+lplRVy80d9rIj5vh3eTLCzR3jvmyQb0/BLXozlWB
SB2sIH0NgzFpF5INA5H3Lex783JRX5ihZALmi3sl4hm65theh2+wuhVOsJNSK/+Q
ti6B8puqplcmVaKUJ9cDihulu5YvA0orb59/IlFAvWwrfNvA6f/MhPQ9UgDE+ofE
jaNbJB/SycPU26R7Y/JW0sRHXmVU59p5aRDJASVMjBwLwG8LN7pwqii8t8D+74gu
Pm+JmJ+D/B8cE4L7lMN7SZGBsMs6Doq1ok+RIF2QFAaEOEmJPzgggis2SH7w/OEW
6jXU9erP6Kzs0+JxamwU3xMXQnezaa7x6H1XuPgiFOCOva0ZA+yJrSE+6FHVxko/
0SOXJoTBy7KFN4gBEiIATCTKtm2Sp51eoWqKWL2k7Lmr5jqggcIjIdYlZ959UzUR
BgYAuZBYIhsDF2ZiqQA55sP5wLJQ31cXJzy63rZV1g7TBK8j/Ouf8twezILNSxbQ
9rbS2RBiJWOaF/KkFFPMA8v72hwuROjbdPfa/EeBtEvCzUziUcI0/0EUWHc5U2J7
jWyuEbu602w3mmy40elAay9mJSpLKcPDB/HUNwwDSsReblDvYlRO3/fud19gMY9X
RGx38YG+A3k2R+P4oJjiyI+xoyJZwnw0dP1lML4kxIOk7XrNtLfmbn9yW1CmgGVf
kfDnEXnq/agGP0U5u6/EOts2v8wjYofHyaQp+9G9IIrBn7TeUnv9mgGvI4AKCDq4
5B6QQpqduLw8akteVI6nMBgKW6Pj2OsF9dnJr7dVK3GZ61iWNT6EL2sxjurOghXG
N0q0HReoSHdZ1kZ7TnQoXtPPE1jSD5NK4c7TIzM2SXQ3Wd6+4JYOFxcxZyW52Yw0
+4Zr7nE5CwD6K86rrr9ZEJ4oqqCqEYby019AvyzFpkwCpixv3rMwLliOyTV6qGms
dKe+Pd3v91BKZ/C1aed5I/2KZkQNS9DLrYP/09KLPUjDs14theth3lN7i3asj5CP
wtwTqdOPyT2AD3rjJv5S409uFA7BrxeNS8Avek8cB++6y+l1mHPt+w9Ey+rZ4MG5
mi4PdwR0BJO0eW1a+juhF6Vjh+/d6uoYhrgIb1qRcIS9bZ6bNRDsY/tPQd7PWENG
wG48mTzFney4paR7It6R/SnHW2tLY9tvj0q9Pkgla8kaETpxPvctxHDWWtgKBaxK
jqPOrVRBZ9VKGf5YZE8SDYtKl9YiVy9f2AnPglbANkBRpSERU+C+3xaLQmCT7Mnf
M72mFig5SRr4W4efK8RqrLbMg3Ugwq9wK30VpyXSF83FaWMWB8Dl4FxiZvLw2+bc
qRFq4I5OwLsryVLJ2Fxd6H3237fN+QMJVEB6+bGX4ku8ENHjbr7hbhf58uhEyhQH
PdyxGQYRcv0gjP8LlHPiQLtd2Jy/SOOgpfM10qFmMduN+486OxG5dWzXlS5fPntu
JEcrdCmazno185hzdqQrUylz8LKLvZJMLmjKJh4n/tXk1Ab4e42lWFW4sJFsBjqD
xGPyOts7tzsW/B1Jj4M6oi6X4FkSNQ5Ev4mzQQtn4aoW5kGCqzlWgVBQY2+YxlLD
lGvh31+8sVAjdJI+TR+/PlJ9F+CWYh/08OWWy7m8b7p5QlGV1YhOaTFaanxy082t
NgZoYeGQa41+DlsHkJK9o6KHP0kaitppVlKWK5laKhb6GF9utwbLMikP1j6c4lr2
iF/rwRUFEsJLiiyUMa5EVRyCxilwlSwkzD3YmA+fsqZMjSOrmS6kjgdYCTHGWPui
R/pxnpVfeZrfemeJXkJL2WTiO7Cvj3Uc3kM/+nmXBqSlw1Z3Z0BTl49vKQKcUvhe
/9lntUVMN3KCPqs95M6TOOe6mWliCsfoNCmE40FB9+598bjG8yS0Sk8m0GviN2/T
v9YwaBD7KZ6vcLZUXWRUKQOXIVILyhAXjh1ZJX/o7/TypaRy7GFHGumoq3PVM818
x6nOAD0HeJswhAsFrOmWL3w2RPGWmeiwGOVYyc51s/2sNzh9wQRW96vEWsqheKnc
0U4sC8Xbdxsi56dramV1hpMY45QsoKH2RZu2o2I+vy2g8XRJeiIo2gpijHwehKHv
W8ntKI3/ZUYb3HTH4RwU3U4y5SNeROmpK1clZWbrDtjBI+r4rBaZbZQxcAVtCxv9
ez7LiszZiLCSQ4elqFy2SaYMdA8ztfm73+NWnYJpbu3CbVOW31XZRHeYJqA/XelG
S3e240k2bEWOueI/h4nWGUU+ugqPORYzDN27M+TRLjpvXynE5LlsKbzoq2LO3mIb
KqPhBMA8s877fZ3bpvngQW7VI/El5LM84ZrXuHwTlRYQhhgaMr3l3ojQxmT3iAXt
1E5GAQ/n9VhDmHWJxGq3npmxTGDRSi3nA8qCyin0udEdXbrqLY6mkf+y6otEc9BW
a1RyX4ZLofckTbviSkSKP+iTcImROLkRbV2OCyQDiVakBC3d71rJrcyUtHtGHgrs
j+5WSswP4ExCiirn3+UAPmqTAzpzaP4at5ZD3VsWNvWyFpdCDP/V/hd2IhoADIxC
onR/F/CSmfBzCXIwFleaulzxuK+fSGZ8kDwaPwOO8pieIUqT40H2/N09sUU/ioKe
C1WAFGNBjK4aPiHc0HHmeAz+Ncqpwu5qYEeZHRyucRrzHF2NFrp92k5wfOCDXjRL
+OWp/ew9CpquxDaxYmxX1lrx7GKEW1fGBaGSFO0boynWySpwGykwPXIKrxdec4dq
62ollnDK0zvOCHzDn+GrBAcLyErJslCUK8h+7t/S5gwjWRusu8CUUn/YkkAKjSlu
2JH1VMF9oVika9eB3fGKSFLejzY5UCmObNrJPqZwxYId4o78mSxxqINO2pfSKoOH
VSjezCiUT0b7xuis07Uvw2S/DVMjIxZv4+COXj2yERgjrolMab6ZHGY64bevSXfq
drWBowgZ6E5AC1vdeF81WFjKT3a7HYkJc9226YcRezip1e94l33qjy+BFqMSqi5M
hHzyjlhWK16HAaN1eNIdc+kdaKY749E/U4vOaxJEA164K+Z/PrRgaPYi0NCyCxYk
sXFbwukOSl2KrdnSOxTNqJ8Xu+B65VMToGGqhw7DamZj5y4dIVtO3DJa+IgL98wm
4C4/rpYoBh3QfmsvtUfZ9VE3QtPvmQ+3NYWxomurVFstenpGRYIimiCwi6AKxaaA
G+eTlHZApr4uNCPvbv+BG3y+swyGKh8yApjzNmDLCUImfnX1ZaOT3EPGXru3K7i/
hrVb4SkFUWMLfuwEsT+q2olijnhE0cqTG13ANaUZP9wYr39VWnfGxxqQZ+XwFi58
SPv2gTqpmj2bm56Mc1USCI0kohtDAwK7clD6eAOVa1urhIZnIcn5laKROwUHOtGC
6uSCDOIl5I0B8mTMjaVEOlvZxj/M8HzPfW4nhsjCqvdqBoKsoNakQexu3R1mLsi4
ZX9TYcBNtQRVESN1R9vH9XrzaAH+RuKhmGHSYQH/TIiooB8WfDNZmpXQiakUgM66
eOp16joL3cWLFaH3kn7vDqJWYqc4HJq3d0+JoAqboVs6vHFR0pTkZgilUxVoRlJ5
Sz4w/R8B6eJpNTddvhJusR+wUs02ry7hr70cAtDP/1G44/TRGaCopXl3nRWfwOVz
ndCtH/Rr8TufN92GuSTC8gmhvnltYKTAq2I7dB1Jn/f7ib6w649fq6b5Ih4Ni4GZ
9sYV/wYHwVEil0sJO/Qy0IUTtSe6QRoRElPa0x/1ukHztvuerOSEErI+qLMTCAQQ
LGWLL9KeyPbPJIwP1cLnsQpyz5es/H7gI7ha1yGuOsMZ2FUVBDICFQrB5Hv8WEU7
XkRW/j3se6Dlf8gaxSrdV3qIm7HYHXYOCpQE862ZDgpf9+tulEERvFuCnrNQO2Ip
gHTWRVnUf6nzRtBt2QqeRls3csjWPa+X1wEias5K/Cx3DlAeI7IHF4Wl61NAn+6L
LM65LLEZoWfr8QWAbO0ezJpgu9+4JaLMjg79+CVazTJt0kzSFGIg8H1cOc3/zsDI
mAKrckf2ETEPN1zwOieBnI4vRWZUgEzignx9v5MrcF+Z4ulrikoSWnewVjNSQrCp
4GOxh2HJ/R1Nvy8/DWil7nlNDyMXsiWcUIBObBinuXNHxP0Jt7XZldardUd+4sJr
0mtPlkh55zXRdjCR0Go1b1VdJJaT13ZyPjkwoM6a3h9qY5hLuocuLGYopvrXIrrE
t0NT4wMYV+EBfpVswjmQtbSx9co7HSw5X16sCU0tmVm4WnUv9LSQ+AQ+aXLORyk9
L5TLDB+27mzZQzQwnGlGUGB6HVtnm/W/M9X9rKRiha+Nu2/aANEibQ8TDa3I6lMa
7rgtMKbRdRePGIpBIr43rcUbsPNe1PycZA5t80+MgZkQlTHgiZ9wcM1P0UfGh4TR
XAWW3v9oWEzR1wbuX5rXRLSVjoZNjqW7DUHH4uPcBckyJcTpPDSEaMBPG6ZDGRfz
CgUsKIOT9DqMOGd+jRYy2hKps6Gi6MK8w30qCfXcSep+BhNwxzoqyHQzyJyroXio
FCORfH16T97tJr1kRIWw8QC1wTQGlVY+lnlM8+eBrbfusggHtH25RJZeEpidxwfA
QOp2LvixWBh0cgYZdvzpcwGrhzT8vlFojNt+xn+ZragAcOCPE5Rpv3xHpGuoxpCO
QPtb+1DsbnsbJfRr0HM87LOZ5ZeStNouyyKQ29LAwpYD4s5KZFOD5ApZtu0tSoon
VhkWkdb65cIvw9+jGnnvi5UVnChtFH5rRpoabSrJUKeXUoD3a/CAbClRNZkuy+/k
1x8AD/x9jKXjA6urY9D4WLfGIgbdeow0a2C87DIx3sjiEdkI/ZsfoqJ4nZ9vn++4
cPGELBkhclfiADY8WK4So836vDgvPxtD9IjsgtrPX+YTBDvkXGe4EXwdkjC/hyZo
fByHZasVCTCaoOqfFpVHN7v13bkDZhAGMjgwdFxF/0lpNGwfOGgT1Q5djHoxuWbt
Y9fEZPoH3CgQVGITKJ1Td7XwY1OkZY19ivDnwDDtaCP9atMkwzLZuvoxAVUMVq/E
DWdtXDTvO/Z3uNoC8GYC0N0GdqMsXuKPDx5wy/OagbLa4+FlNBIiVeQM3auFAJUX
fvdr74X6ms7dk6XUwbj1dqQfhrrnolxnnTd03aixiXNT89ykF5Lv1F7YFqnuo4Wg
GRINbXH2XZAw5xVatcSjyiuQ3XIAQsO5pJ6/2Pr7zZm3Ej8+mKLmqnaxOhqRxWyU
jjdwZdoDixfij2avCtIO+x35bn+SRcn6ow+hRY+voUDubcUF9MTz2ew+2ZCUuqVn
yL7Mh/ih325fHDCM5jMnhLDKDHO6v+UB0T2tt9zFG/JY5f4lnFYy0mr02esSEw6m
U5L6gLmphldwYsXDVeA4bEdKgisRa1aH9BUSet1a2E5/SMDmzm2BXIMxdRR+Cxte
zuGDEbiJx6ryH1pz4ySsEtwMr2+3NAa3xLLiPMm/B7wx7jZu5IX5WsxKaDg6chZS
GvoR63UTNH/xCzjlW+1b8ipjhjvo7zUQuomDkdM09GqGNhqkzkH6tNXXC8Xwkv7g
vg3ZtsGIKLTVyG6Jc1VbBby8kd7oZ0BIwZS1vZFBJiyyvTOJulC0iOIP3KyTgevA
P0Rz1/tWvTo59jquYz+vyYe5iT9qM0YHCx+MNJ6V8iFAthTY5G0364GaiOFW6U2E
LT4L5EsCrdkffTeu8lRzumvzt7gj8sOCSSZgTZEWPgX05mbpQeUn4XEKn/mFJSAH
Tsz8A+OLvwe6k2nboRZksBfyvnpccFwarJhMXlr3yPx/q6eROZceEDYwpZetwoGe
S8N531P1+yuYNCP+QX7dkqlHOdXJJyniH7h6as8fzRQxHq6+OE0KyMyn0W7A5S5j
/O4l9xONiZXOn6cLlJOMV/tBY0NMTsStL2GoOqyz3MoAG5zSkYLNjxiZpGApVWzh
IYyy4pE9aL3Qy5Ub5t3kGmTeF2TOSXcPfFiw9qAmZ/cyG+Jqv/Q4QLFgazciyM10
hNCNOSvl/gNAAXpt7G8syp//1dqdxFbiUOmN7lLsWOl8NIWJ75RgTBGp6yPQUFxI
kO2+OP+OHjgK7ARp5FNDoCXiSgrMUSaqM/cZ5Rp7ba3KhDYBnUteiltTwaUOvJ4n
1pw51w2fyvgiScazpJEp6MGB8y4ScUicTTJZ65lDEAK3xhy9VIvEVj5HLaCbh/Ha
R7Ixurf6Gxs7OunhxkgK8wYesnPfC4+ThUwJw+0kYrHNyoRaGGexf5Z1avn7D5+E
69P4Y1x4nxysLesiThX4wgc1ix3dQZ8BLaNsNnheNMrfhphcpqGznKOA3tkshHus
FHAMR3GOMjfjQaF1DZ/Uf6aTY+iWwW10NiFqV0hDCTnY5gn5l5vghtOJSmHkTDYl
yA4FFy0Iqh1cUab3xJ1FRHt6ra02p7zXZhCN3pgWsU60PP4/6RQG4MdLw0rxsVtm
gqcXC12wSxJRciIv50d7P6+6FmLs6RqRdH7weiShIMkLWGVRytbrgzBCHoeuqwiv
44EjTtVzpcDE07tw/wn2sz0wsQcW+Beg+TzT9tXRq1tQnXXYJoWU2L9FkJUY8bnU
M7QIxQPWLW3otum92GS0/Tx7OPOAz4LHNJmC9WK58VIOhzXUUEXdtqXKXO3r1+WO
3cGy0NOZp4jJXLXHDHld+dMBcdsif3BqSKDWgh5WpR8tkReIsX/ZuYa02irQrNEM
JsgVe8NQp/5seEJ3+hMZjWWY3qUrK2621gc8xdrc6gM3uPRlYuUNZ3Gkt1YF/zvh
TybGY/jkoIbusgsK89uhCTo5pYEs5AaQd2kphUIzyTihnJhYiB9ucMCB5yjZTURL
Eoa8g0az+eqpv3GtIwUmU/V1FuJwfIeMvDq1Se7mGVxADIm7fgkC7bxD/QRw7eGX
0Ogdb86Z/7lVioSh+Xgr6ekmaof7CvcXMCzl0zZA5YY1j55kktbNfW65MBrGAmAc
tP3mECIcIQPqbRbp3O6HPkLbmpyfjfoneo/jxoD2Su3jBqyAkzE0UxRp4PgDXjyj
NvBIJEjdnTgvZu4RUO34L+dAWp3FlupTtafenw+4I6VDoFCz3SHAjZJb0DuVn8HF
yLqFt+00jTIPy859pdva8+ghfhPGhim+8BWD+vurSK9uBFDFvl7iGyc3xdQeOhFi
mKTpvekyqbSDlRclawEJ6IphKkzeIfOhdzUrn1I2Y98Nu4SLut41N0Gfk8oy4lOQ
Moy/OC5abeg66OveFywHyE+/hVg/OV2LwhTxAemSxcBfTGYb9PLYfDi9YbQenUcv
OBtCFrQrLBiP2rn+HfosY1cDP2AOn1/+C8IuZlOY6ymhoRIkdpZ+apGrm7AVJpd+
wwfbn5LRLxw4BbGFpf0zNrpuPpbj/yRG3MXAnn3lJUzqnmw2zqxFqajIpjn1PMtY
E7YePCzkzK7vAf4AtK78N/tYBv8l4pVmI0qFDKma6VhT+e/zZfcjwWl6e0nnvl7a
tVkYgULCbEvjmRs6nQvwHp/ewsJXhW72jPKknc2RKvsOmU21+7Lgh93pzB2KnOAZ
rJAg2swaPWa2xSNUeY+fUWn2TVQy7IzuVaSrgR8HYKwdBEPQoka1ZGnX+QBqUxqq
JoZFFkG3atdSciJ+Y2kMRJENatPBdpM1adzdbJoKryqdi+dTC8hxOwGyxvXorAp3
+/b5++jvPqk9cMlvRNAbT6c1erUiMelKgtmdDJZXjDz48HN4n6R+5Ba4J+99d79n
tE3xaaSLhwRuaRg0m+L4I6THfQa8vR94QsInYHjSrvL3bv1Nc3vjlBBCILPiJh4u
aMQTYROtSkkAho9dwaIcGX2WgBe5XDuvnYR8wNSNaURxzY1owIdcKAvlIUPgoY05
fH+WML+eSkf2d9RC0gf/G+0oC27iZ6Sd18TxRP1ToOcb0BKAjA4GYqwEJX6MD0Eb
0+AF8G0ZWtn26Yg+sRyd//4ut916jr5MuCK5rWOHLDPfd7cAwkk8k4G8csoXsCaQ
3Dq/yAEjFUpkjQn8XoXBtEZ6SLYZBRDc+zjDU7h6c57H2KKu+hTNRI5aZN2xsuso
0XTy/pXnpUexsBBJK/iMuY2/cAQfdFqwhtrmw7S65+8DB5YP6voo7nZFmMkjn3BH
oOYMSHtl8mPXQPCacCTo7bcCr8LKlAWKeCiFrYpm0W0znKoIyXnPanaB1jrh9Mti
Ds+Hz/TRqGnuT/JrJhEWMocy6epfdZawqa10EBz+poKoRzdAuthXrom2PyhByNvf
0F5pIiAGxMdHaMltYYNspcxoHWPQWSGiMFZ4whLUxYYjCRJq62sAFNJ0lk/oE0BQ
IOn3GgZvLo1BK84JIzBaPk+t07jLkzbNRGA1Ns4Kxpj19v/ply02Ayl8Mf4BeShg
cw7uDtvfz3ldZhiuL79IrRBvA4qxQH6uEA8ouhi2u0hG/KKzD3ml4R8JpN6zwmzZ
peoZH36fbdyTfm8N3mtyCYTSgMVkeTm17wWscgSwsT4ydC8bNjKyzRGA+aBXm7q8
qb+lE+L6yHSaPxPIukcBdmJ7sQTMC5u+R+ne8SBuTX5Bf7dmgP0MrXfOPzNdxadr
GKrfmgoVC+6rrcf7F+aldXYkEFc/f4+7Eyqiavd8fqlVDU2qJwSxYHHqVue4voqC
0bs33rp8jjs6XdjR5rmM0tyqiRn/YXLm8KWid3iASlaBacn1sHOG6fCvByj1xvUz
AYWK87edIFsLCBjOjLwprcheJ7WA/pXhkiciSjemmWr8kpHGjlsh4z7yZ6URgA4d
iu4QTDBedUcR6BFyzr2Df86Ol7hqaPeUhNW0A9m356roKHFUqHIFcmnFMkjmpysM
2JPTyHbBfg0LTJGhFuQg5Z9FtxV+L9zs0rqxtY2X977MoWBR68lF9fmhodWxQ8E6
kFCYNTGXGRbCMQ9Pl9FODbDg8/wY5flZwuH9mX63Yea2WKQpqVeZVYNQXoTeYEns
vRIcs2inUXVbBR6bf4o/E31Uo03xjrLm30s+Gx1matvQEWbyNg0yU+tdjS3RdsZQ
URY6evv+RUGLaopRJsyhJSVu/L+51mq8rvF/AB5CaLzvBIrmQCna/m82QAaYLizg
OlYSE4tkUHMvWdPPqD4gdgE6Ycmj8YPLW4Nfl5ppZYPh2zymSFHkEPPusdy+cjWq
3pwCmOEk9xagHCgURtwLCSJtKSytJhe3pZJ51nXXdQ0vKnsN8KOVXyBX5LUNJy2p
dqI0VxQ9o1ObPDdbN83jwqIHb7NDVjMaH1/utPbwOTaVd7XLJuo5Fr9qaiJd3BCS
UcYFOg7k4uluU2rboWgsDUuLpOtPyxZUg5WnpDX/3k8hrf0wY3i2inhTEajroXTT
VOUYUHtSN1PpwQaMrTX5mHTbzRr5/27ifuFX6bfQvTpWu0jSWI9bp8m30/G53x75
QFnliOvk5nmrde4GiGsoc7H41Z5oAyTsy9IWT2UKcOp+4xTUDdXBY6/GPCVNQOrX
T9e0v4peyWyEm5O6wdxtVondaRER4aJNc+9pI8dLg7Xc5QOBe/SwWuarFXblOvPW
TGzYuDMfIEJl2jnZfoepZg5WKRSv6f5bGOiX6QZ1nkH6LssoSZlkeQYxAOgTCOJf
Y3gLKPmyQyYbIAVkZJFnqx1X9bKwDHnCpHlsuT6UhP9znf2pHR1ISPOd6V0BFhJE
2uzykLeMqaBjvNAjbiB97rrGLnw74qmzqwKuMtPdgqMFtgRFYhGD/wI6f8o0J0pI
olpiQjO1E4EgAV8ekohw0HYAc4QAvdiz5AbYJG8gNeJqItbbzErk31TgU1xq5yCa
AQ0OY2sV1F0PRfI9rBLS64asBZxNlRzHvPzYvxHUiaoJomWVCQfriNE0Q/StE9/t
bY/qhRVT/hUeD7oHW2omrVNUtOe2rxhkLepC4IaqZrVDm2PTvqu6vtFfyEACZTWC
/IxIen9Xpus5ZBc0LlCzij5rsaeoXmjJrgFmQXjto/1NVn5nWI5jO0ixHiGxkl0h
inL+30nuGL01WqD3D3pL/FnEFgOYlmciW7baCxKqJfofUc4nHydI8np+dn23jGwZ
J5JMJvC+UObVPpqDUaGHkjU2MnMByC42+PuaV/RgvJn41Cp23p/rDdne34i2tW15
WTpJPERhi8kAjqF9eCdaaEHGn/I6G5K77t/CLPoBHdX9GJFpo/BeVZhw2UXrsCSP
q+NPPb4L/wsRxSryAJes5lnR102A8L9XExmQh3GyK0QEiJ154W2n89RL3VfjO9+t
aFc/EsNbsdlWCbBc6TK8+4BlOpHzxqpfu3nXe+rnfDXNK+zhUCE17rmf/qpu20+d
Of0sbP1RT/dvlv1sSND0iJq8jqJ2AToR0exCmwaU3CMyfP+8KN+pgKqf+h/3UD0V
NXQaSARpTDYTcINejESAhKgJUcyGCPROcd9Ss6C8GypP+GQ8mQyGIunXI0zC+JAw
aYf58XIfQfCZhJ8zj5r/ll8CkdJdG96gJp4W93PwgNf68np5ZNpIzsyGGIynxBDI
W7iEIjUXFvYqNwAWsJUVxiHFkjMhxq8JtlycSedvaDSvBl7R9zo12kfn/zs+Q2eQ
giimKsuyz/WMwk7G6ADpPLnJrlnvDyY5+1rUi81idzAIX+ZRi5VgrmSAu/LbGt1x
12PwtCAAMWLODCZR8V98Fyat15VLfffj372IiZ8Bc6TgH7yRrxODSMRkSVn6bf+8
L0X8LxwNv37jcFq58UrzIzaygi9gmSyoF1pp4cMJGgaVF5T1lqkkxaKdeSM4dYb+
vHFWpZpZFjANpPTGfY4QMXetvcxQAs6OU0ESwFSTD2sawWOPhLsIW/ci5o15BtVu
7TwQTtjmEdvwfkUdvB65lOupSSwTUZAtUmCqVXwQ6m10CPo40of07Msp8hm9YJLK
tUNCC7FQ5LxxmYMuODw5np7zBKnTiforRHrmmNc30oM0rpbBUb1kOk2RCw36RBRZ
FPsajD52lFZmComAybdG9Feum9SbYGfrx+esKYM6eXgM5jhsmogQ6/hN0WSfI+lX
s6rcINXzH/2Ol1Ucgydf2NgSHoPJP5biaizoj0uxFQ50EhgWTpgnOErDqrFzkuxR
4IT+43vJckWHKYjFaQHSduzbB47eGi9hCwYokfIoMp1btN0vGNGYS3qZfxFZXyRk
+kOhXU2v0ejBPUHVSymoHXgRlajugw+h58UW9IP8CCNa7FHC3Vmet4T+nsGx4fpB
5NXEtgDEBjxCUef7Dyvs2ZMXTsyur/lDa1za/GSg6u0khNmk7HDskWPf4o14fn0C
FR3Qp/rspLDv0x+Ep3fJDt4vGuQCLQYzrymus6piNWCR+x/CEEv6q+RLaUD6WJ14
XVatyq4xitgVIv0HZxj3asXyJ1yBSTQhd9FnU58yr0swL9UfGDF6AnkUMKtLlZyB
soOX55Tl0sF5aDTO+tTy2/XwbOdX+NH5QuXoCWhm+uAJLOf4xZDbkLBZW0syi4zZ
LMMz5YxGCVoC4ZKOUqlgO+wwnYGhjP8aORzuQIMKMRbVk9Smn7FNFVVKodeJxbC3
g7QAI6IMNE6E85z2BtluBtU7KxCkfA/WxQ0MWUdE3wec5pQE/iZ4YkOugIMAMFlw
1hlGoFLAFHNUYLpZVvLw8qY//sUywYP11+tLfdhNDQKXnvsRKnsINDNAqSzJzBke
nZR8iADZGMOX2OnsZ0MIb+ckaXknoEW5b3O+U/SZkQnjsKKqNSlAujlRRI9irHUC
qBWzmoWNVDdCOG3uKmVmIkf7EfmQvSFo9wa8YgDh/Os10xAWy53N13CPtUYioLDv
Dx6VR7UNrYnrlkY2Ne2wHgunB8j7eJL3aOni8U0y3+G6Xzp1QYIqdF3xNaxC0L81
0jxy8PycjHKvGIfi4MeK9V39xmJ3GKqyPMd4yZA1vyKsGV0rIhR1ZyA6YlMnNPQV
1Xf6evwtBGUerjNqA2EL36bjYHvV0ZVffSguJzLoyUIgOn6oeIB09YImdo3okIw8
Xdh17lzsKIqNJ0OGq97h1tGA/oIwJf4fH4i4wfYapmkvjQzsm+2plnaHlH+wiiCD
Fpa2wu/SUHzWKIZFaHOcxwCnA+A9Wf1sp+sh4l/eGFr5DQ0aARHSECsOEyMg5Sjn
S1N2qLMF670rwtxCq6cBTpfYyhc6o+z93FxGUEDmxeik5xSzWI8SjTwtEmAViSTP
sS3ESQb/L9k1YuUuJ4ou8Lfy+RvtYPADZtn2hvNG1Amm/nEl2ddi9+izYVJUqgPi
qsSdCfByKOhP89PXtggyYLwN73uFgMMPeFXsCaKt7BgNTCewWFnCjtHF8Jc2RrXK
G6t+gT+loT0lALqOnyTUT2/8uGKmCt6wIhWW08a8X4VZiFNrDHpj+USgNVmRCC41
HnX3N8kfQHwVL5d3r68XHTN+uPQUGObm7H9+KHGoUH5ruT8oXggEtGGD82XAPx9O
2qjEgIObCyMLbT4xRW2g0D6a367WLdr49ahn3gf330c01gQHfLuBnYyJwB101RJF
jgjM762ZnUP1IcaWQGj3XR6aoYb2YLjCOt8CWKPgci+Yz6YBFmpnI2UvqqhjFaZ5
j0xLCgbqZkcb5kBziGHRZRSpY0y008yJyQ3d/0JJPzSTTc20LjWh0WrZ7fjPUsdF
Rp0Af5NNL0O0TwAkRX8vKUwMBmYO4ZDwmKGBwFlxgBsDGxOSX6BCaLGBRd4/SBga
X/dJpnwaM4TmiHvq67g/KiO7UP5FXp9P5agYCL/YQsPB++o2sL6WgkiHG6Cz7rGL
1g4adn4GRCg4m00bIBhRKSfe0/1mz8H6zs0UbT6iAUjrHiESeIEQi2uXKhbna2si
DCcaFOvD8jYCYtkN6gDfmyal5jlZd65kj6kZEZ3OE7JpwHevTjrV6Mp/023lZost
gsoBqCTS6fLAA5/I+rfLzZl/ENbeWq+AEw7V+AcOVJTwC8ZJVLGsJ4kw46t4BwsJ
OLgyPHWU8sjd7Lv6b26/80/CF+AByDsyqLpWH513PAVzAcAjW2gfwf+FDqDzVERV
3YczN6MoORw6nEb7ypfo9pw/VZZGh+dVSq5r3K5uL8nDnTtCSRcfXTaRNlW46h2n
zE/tGR9e2ouvL/mrNjbl9DdgTRblCOMF8n2QUcPUyI4u0ySz+NToOa1Wb2U20JqU
Yvoyv57VsKjmh8YoNoyT364FTfK/6NaQ2KJbZV0tIJ/cj7AdEfjxCtpDNk7yInI7
+TgBGnJAMi3dbxhsnryOx34i0HHzJSPmDEDX9TvpfyNFtb9gCjf2vAEZkXI7VQEX
FJoB6RPYnYEISEVmuephwljNsv/rc8WzsPdKnPr9rjrwY+qu+54hRP0+d6m8cwTC
YWyeij7TegfCR/s3YYhtL31a3bpWXhgKulxny3xEQY0MZcYkoREj+FDqyaeArnDA
UakqWBIdNLPTPNdTx6iRMy9vgR6wIXPD+C6OoKvU3MYFdImr/C4mEy7s/UFCw4fd
39oj8qSKtTLx4P1v6loAl8Ol8E4raAePBuvDDZAwajFjfhgIU32qRc/qmsM5QDtS
gMybMvIlbw37hFe96/n/TlwLbnQUmvX8MR2Yq0TdZ/FEOcqul2ar9LsH+eESm9tt
RKVcJCXqR7Rvo0sSIlIxpyV9DKqGiknkcD2vPCGNpOdOA8rsqn4d7rhj5QhqizWC
cytqaqaJ4W/TrZBE+K8nDYPeKsoRYVGZGPzl2OmbrSXe9OiTA31pSL+klZLcILts
mehy9NOudEIYT6ZB2iTkwkEG9S+NbpTywM9ipxxQJP8WMiBlO756DBE2/J+s21rj
WT7ETlKuAvYcZhlIWWxz/wa7VaDQTHL87YGTeakA/gCnYnFT7AIN3YlJcKb2ipmK
gH//5wb4FbgvN4uzLomlvmZekk+zursWohNwju+NnWqS82DQ4gP4YleX7WcqOGtW
c1PopWwEOBU4uLd/gCopS3BhAH0175vwIcqK+niKSJCjWNHMR95nRpyyS1RuWSs1
xDt1Ydoo64N/6l+bRYKIuMoE6QzyLpJsOVd684MNLvB4VavpAcmi2PP5tKV4Mpj1
pKyTQih8JaKX859jvYtbPCo5aKjsIgyFVPNp9SmsiF5zuCy+vHxQefR9tKgvk1Kb
Ml2fJ89NnpvOV1byb9pBv2Gh80RxyURMcTkTMx2O6IpfFKax0A3FjXdHXXLAzgyy
2c/fZ/KPCc7ootpQYMgIAq5Ah8RJUJbvQmusaXWCMdOK0lsXxHT1uCFiLIxGRrje
kbyZhGusCRxHHjA/rAEMmoxHTVtqLnjzXrORO0HMtCAXUHzgQg7uYrSTAo+b7PEK
JZhDpNZzr+1ypZwbMT0XpEDhymAD5DLq+EVqdtM0U/UN5WapYfhIKpkioo+YAQJ6
vYuCwZFZ1wo1ko1jBYMHu0uugsVdhI4+ZWt6rccu8WqPuBOMyOGeKWIpMT41xPEu
/JJa+IjmOBFIO4snf20/NP604DABlhfiJep/109D3nc41QMu00m+UTg/fKgZssDA
xegojsrFmIdkucImLuFycfdH6Ja0N9q/TaZaPWWGpY5o/Rz+sXp6b/+Fu8xP5vAC
2iJAKo+eCAL9791EY/EKA0N4+MAEeN6wobnuXVwguQZkIZEwH/iSnkLDE/dP3oK2
Q193CsFVWyR4eIdWakZnJRhLkE7mfM9gssDW2erJrmZn3z+4PYN8gH1hMSbc1NLs
6nVTQkWZBt6x9O63DT9CYMc0Tr+GIqZopadfRy4j+D3Vyc1p0LEWztWEOvqTKCMS
QhrJfRnf07ka7PmIeqtYYAm1RySafFUefAti0/jyVYBj3y6dTgojX1s3oZ7C0W1o
IwEySQp2bboMv5qpLuQEsT47cqB+gQoeB9sKUNyIJDAuCxN+vnhXWHKLOgL1R+vP
PIwi0h32BehxzLo+fI+idaZCGPo6YU5TckBWhAFk6+nSaBmEWVOgxukTlQ35qyyh
QmNgHL4iXt457EFllNbj6N5sYbi4wXa6+/H4mrHC/WrXcPPi+HjvwNWOWaFKqMoe
VCe04iRNFt14D8dVUayZ7o3NDY+w01isirlBxsLrX2Zj4Cs/SGACPv3gaYakhMF7
kJPPmoOz7foow1tFK84PAXYiDaOkaB8nguXZ+TlC7vo0Ba32M/WUouSDYkMN/oNL
/i+BkknM+X2SyqAYbbGglyKnR7AalJRdySAMYc7E2sPcMa07wqA2MBN1N9dGs08F
0UwO52T/mjtfRe78GDwofb10+tQEOhdMkVz50/xfaGxmgl0CiDqY8tWZ4iNoQOgy
gg0iaiMdR/v/ztVKolhrFGj8NpYfuhSteXMxn165/wuHyWUR1/LZCPpgDPwCsuow
+MxoXmmeP1LN8cYqe+M/lGJWGpdF4LSzrDYViA1rnMVdMRvxQqo3rpaeFzUDrpN7
UyYucKcmje60zo6iYvIvRhdc5Ld4I3ZNnK5RhfnhUxdt92oYSABrkicqoPV6+yOn
AlzESaYNwhW4wrnwZFsSh3I7RASzlX5iWY656KWkDDfLoLff37q8xJkME6o4Cobb
k7OlFZWM/qD8A35PFChgk9aRxXv0bV7J1uddz0wLDI7vgD7zr5TpRe6sGrFCN9Fc
7BByFavDRG1RrQzni4DepyJZMN9zq/UsxbYp65YLtZzRuytR25zG1BeTRWOGEopT
DhJ+pvwi/NZh4r1eovBxKTE5W64ZVxmlx/ojOntwEVt/r2wDjV35G2u1e4IDXEiK
JhKLa5/ixxJ0KKEfRJnAJ583QNtksOFe0h4303y+nSZFc+CXxohAqHlnzNPXa4LO
VVeGGqQZb8+fNgA1/KveKtIJnENzUJNEZA7hZ2zfIvBWu1fk4MP+zJndZ5mAnsJ9
CWsMROknwH6pJnkx6jbSOqrONm1BQeo1MJVxP7g2NEuVcQR8xJ71tF8e9wXYlGq/
J/LfYmiAbBAjcjZCscFqWQayAiZ69nthIMWI0SSoR8aCkVyTrRBwtn4dLThSM8f0
HqZScMGgKnC6qbdmdDMp5HSj8akxsKSZLbcmpHWOMnWBhBZjwuAnk0kHKS36+n11
eq2itaMT3iZJfQ99mpp3Bb+bwzB48d75z0faA9JuA1pyEzLM+7LomIZRYcOU9cVT
Bdk1JhPtev7TvcFbiMjUmZxtrwmm7rcaUOjoWGK0C6HddBQgbG2U1XV4ymOQ4YBM
qUrSI5VGdm7GpXuZibIEichWYaZs2q/8hDkmqSC89PagczRbr0PaNC5cnnBQ5BdV
52Qvobhd/lGAvmBkiL8bXuH5by4tiG8P3ESZhPu5NF4WtwTXy5L7oi6+QTspd4zo
jHra8HHbF83+V0If4i4Bca8xBHXABCqRHS2phzUa/CsaXTcid+ijiv15xvAn/8Es
EuB1jEHsO6674WfeDjpEqX2APE0NZdkYukWJxcWkDA1iGzTPo2uhckxWrn+e6vwc
bOIoD1ppmwVjXYyIqiIT+geel66YbLm6dXY4uAAVsJJZp8vphElBRjQqBUlt+2I0
udl1u2Hj93Z/wQZCMaS79sdRJ7Sq7ZS9oxMWrZXMRJXckFQriE5+17rbRUzieeRr
gU8EdbVUK/4mGJUqgyPJtpxIzqpw89HV/tkwlE70Uax06MJd2t5NlHQizEFguDm5
ZjpcJuRyzD+pAfiE/eva6kL+8mbt8q5FvgYvaATujzv2Ntr4fvJ2HvOGnB+OkgnL
B4O6I1GTVXx3SiAogPrZYK2Uu3wSX0g+ihHR5v2A2vmZGa65rrePKgHTJvFa2+u/
eIo+adjcb91e8gADNJ5cMKc6+z67WJRAmejApQvr4tF86uupx+IKp/IL8Gk/T015
589NkZVgc2M5XYwOXqyluY1+BuoMWCqqtl3+ICUDCaS8kdQERVF7Zadye5UCZ8v2
hX1iE8iqEOAdSf+b99megB3PfiKVN3+VUMRJ3uo6ZjXPbnq1qRbDXWSyiOSErP8N
PleaAeCyawJWCyeROQyv/NsHLk/d2++W5lsqsuNvsmjZJY0vlxP6o6oEDZ8vPOuG
wHpt/9JKLKVK5rbSQqB68AV9Fy2v0kRLITdYaklhuBFXRNm5zk5br7yk/EkAxZQp
mDt5EhisuzlBycuUBRihNrweco5u4+w8WIKJsY/7hfPY7jUsO6p0ai14SGhe+P4p
5jq8E8ku9dVbyRoL4B/kFYS002+AaF6tLcp7wajTlqsomSzJ2pn7noodMELOVeNS
pFobgzGcreGgycD74K1d6geDy7sXtj8lKUs3JJq91nYnhMg8laNdN0O5OVyY+esa
InOtBY3QzbRZVYf2FtF+fYwzptarxzHbCvi4aE+5XGPM4PIoscUfh6LRwArf3vx3
ghCK/qzG8gPRxLtyMULNSVshoiHvnA5qPnE4bBL+K4hMomAptDXucpvh7apwaS69
pN5EhALf/IgZAiFDzNO/RTx2tVjnmnmariTUGxNhHMEbImldA0QnoAKVf4/pY9gS
O6gmL4+PHUnufZSNlJ1twkTPEbUPg0css+UfAieAQ/9mOqfJDSaNx8KhK4HITXv8
cNsLygVR8J8bJ8227DYA/ZG4W5q3xaYeMq8ieMFz0W2CyD3XvOfirE2iQJHL0Rif
FmmqlVw4D4d5vK8xzUY9luk3jW08CbYM2RuJNqT1ZpqFBxDRRK/k2KiiO2Z/iydw
K81jB/Q9jfN8U1SDywSzxHyGgLED0dK+9l9Wkx6vvoAQQU0NiFvrZXsncsfPrB8P
WyoYKaDCeU+vVpdiPFcckiNe8GQxIaDqtmhN1l77f4qn2vTHIS0PS5Ol7nRLqvMx
4Z/BNC6hIbX1m/sf32sA696X15UaOtisZXumjcRH5/SKwhPdfQ8z4B6CD6v24Gok
Wz4tDVuaao8dA9xxnum7xVtZvB5NJPeTXlov/0+wSphd8Y8U4ukAJuZaSnlt4aB1
qARCJ2RMOhNAx7RR6eayIEl6CZqwzCL06wZUOiKYFRpb3VlfaojnGz9YFlYZFGYu
rXTK36XFnpsPsClXi5KQTrMOFJBoeF6MudJj8e8Et3XLVU2c4zzt73ebReo0RgdZ
vNJl5LL4lvA48Bm8aqbktkzTSyImYEtovhxShhFZqdtcP3iPTmHyeAfYu0qEZJAu
PDOWTuybQ2L6tdoIiHxcaCA4lT5nQGXonuYUdQn/T+IyDdzHUXEbMZEOnwul7Pyt
a3Hnt4TpMxOIjL72Pq5u3lf2stoasaDMY1WAkXX8Ruj5qyqNIdYkqlmnZ9HROjIR
uNu3o20aHmcBzHqNLMdfSocxvy+qsK/FECtETv7wJWtVHoH8nk8BR9Ej6lKDCfoW
pPLQsD0eKfQMKuBbCm2opiji7p2ndszFSh2E6JIiusJPf5oImGYpfVJTX+OL6MvO
gkLea9Nyk+ZqyqogdcVOgDAiKYyuocSYmXm1iMpUC+lztZpTBSdRHrhLyCGcqQGn
+bqvzoikRL7KqZuMsZxwW5MTj8haxHA6m4Z9grJv0fEL31ZnvXP+U5cxGHkysKKJ
MqAMX0NfRdDe7nDPfwdsnAgRRYeEfXuTSv8CKpKDF7tYljeYskxpIKTzBvNPk9ko
vVl4KvW6ODBq7rXn4scz59BlhAue45UOMSaA8r22NkflqaE+fSofVahHWn4IB899
9RdXQ5hbjq1reoJznG4/GXXmv4Ffkf22+x/uaij1N+5UgOrPH6FcO53gDI9hZ/vD
AWXhLOP/TaGK999NUzYopPedG4XYZhAueU7ca7XO/YjV1pcPkIZ06ZnfPPpSqjyI
ftd+8Ruh2yd5OtYOQulql+UklqemOSTO2H4rqIzEAkOSuYNamb87TlJ49FhmaubN
3jhXZRrXXFIRzg0fczKtuagrYJ9ZYQjh6XhLeuvzbQcfb+D4Qc/q1Edfkh2i6qNW
oJbxLwJDvh4Ya4atBhNng3jUMpamL3zoHiMuMp7iXpryUHifa2lIMAbN5HXbvclR
efcslN22Mqf/BYKselu3AUcINHoo82rilZneLrsiqvo1RMwxCwvsgMSKVgsuy8Ic
L9gnV69oVebLd5GK2Nd792q3Wa6UZxgTCwfgZjxYHMLGVfxoG47xiA7dReCpTNFJ
UQAEf9D7/NrbaPYNcs2B10mHtId0LVr7vcNiYGCxn+3r9q6LB6tV7yZTLQAh2Yfv
MTz2+qam3Y07EZVPb4BVSUl6+yBQxOfzD0WzwO9wusjfWQ8YUaarrBSA10d1uNIm
7Zv49j6ZTo2eAP6xKeWOyD42fEl5J8s5ZGvgZeaTuw7Ok+mY/LtIpI9lN5l9FUEv
MK7I/OT3P++RjpvEIyjt86UisnGP/4qFPIVo8tMvVqkhbSALTJ20hYvUIubNkiM8
g1HUOVN/Lntbort7uoWb/4jQyYaRkNU0kWZH6x6/F/pknRiKYRRmO9enK5DwMA0K
umkKL00HRisLKs6mdp/ZP+cRwFGibsFp3eXq6H4i7qKLIq7G5GHo8IscqLoIWcC5
7vCMwQ/jQ8+iKo6T4meCQksUz5N00d2cMFfOBDOGGJbJ1TzDykn9ptsQTPerhkd4
l8bd5LyLOaVYCUBRi7pxF1FZtcAM3FPv88X/+05otFUPlTOKeX3O5aVKiwUrq5gB
G5+iv55btyTCHlMHyGn8JFfpIEGZQ4E0i2hWga6nlKSo5IfEsWYK+GCssjtAX2vn
r9Spud+8JRV9tcOhDvc7pvoJU+MkSXDh3NnwDhJ851fCYWBcqDdhyZ1qM4NRGoDL
bonMJv8sGEqLTy9Mp1xG+LX2i6MuB1S/4bXvWxiFscdXYFhpT1YXr4KuZhD4lZ/U
SswDZt30ZiDmOgodd1nFhLVh0vWHbtuQdQwyxh78InNuYnWnbgIyt99Uf3zRYbGB
VRtisEoIe3oGx3z6ErlmLLqHNOIy9kR+3SBNv/gOq8DLeypkOT/C5VIOkmIgr3vB
O/5s7zhVNKMFx33Gkb5F45H9KYNxN6mpm4c83X3FP36ovUEHx4uqbWDT0AhpXErH
fcLTWmzJ3HMimQg1am//0FUp4kuZ+hOlSppRaaYxKs44RPdtJvmbepqYsHgpXxkK
gScBYlconGYrWf86WFaBybn6RgXkO73FjyQ6o/vR102dwKCDO2H+JtN0Ow02xif7
SYFeNyNSj3WGHQYeslMBwr6H9Uvvbb1umFCYaGK0Ib/NpTpzotVd72iQgKW3Al2k
f75n4DD+eJ+06v33gI43+LtLpK2Au8O9oBvlKnkwOKmEeGPHqoUyOjJjxh+bAez1
8rlcquy5hx08ERtkvqxXcS2hWHyKJw97m4HE2dR8MUkOZPdLWuzMPbM7jMHXApbX
b+ViH7rRQhKC+bgPpmuCinCFs9+PT1tVJVM+4wwPNzDBMwEmnnRgKbwUvl9znx6o
4QgZuqWDLhu+u0MhGBNFJKG+XX1Qiujs3mM9Wp1SyLZYC7nPL2K2v67uAGQE/CEu
kQAzm+qvtyDPtYvaNGdjSI4pdMRIyycc8QPBFfpGkyvrdQekRMLLigPcEnOb7WP6
gohrEif7kpOH9MbJRpzWnbdeYDj8ZtFDJLSKkzbIhOYwiPG/z92kDUT1ZDkV8lTX
40jPtWe5hHvMiqfY7AKADqSfN2A77X+gN1ojBVDLuvVb2Ps6cc0U2kkrBfuxEX0/
zO5CMM6j5nvYoc6C+20+4za+4jIZrLxHngIK1ZW3MWPARUg4J3mhZfAa1KWHxksV
zcmN86prudVztkIVcZqz73rtY/ohlFP39LhbT3JQIhOu1iB5JxR6x+TmZcY2v9Fk
gcGTMd9n+G+wtPlkrM0OheobIP5XEeYB5NIPY9aysQ6toxw8OomHG+AAgZd3cILR
JFhY/LYK7V7ehDWIyPSRkwZcAEcMqIwyD+fjMjWxCC1136TFdF0iXb22Kci96TvX
UF58BecOPRC8d6Wzq4IplhArfEHMWIydmqmur9u9O9FZ/Ay5qkPG1U9SQ0WcVkyp
sM1llV3+ql4KtRkNsOeiaQ==
`protect end_protected
