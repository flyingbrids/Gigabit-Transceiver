`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Q42bN9XXpai+nNuVTAcDbBeqs/oTIf7HL8BdV4bwrDtvv4+plSvKkoTySetk7gPR
VpoCo/a4xUAng/zDF2kCK6ci6uL08mJE7L5T0a6oqi26Untxab5pB61j/xN5pNmS
tNZ+GwgJZQyC6eHVLePlmjTFcSY6nSGM+2FHHdWOfY1H9Vq5P6iYU5pUkLY79ma6
NFw80MTT1zY4mMm9t6dPR3yVSloKc35Foc7f6Wc8lr47hWvV94zw02LFuONvIhjw
C6D87XvSO0RPiCRIerdAM1sJHUyDSoEIFTimQB0RFGg10HuhQXDDKv+PGocbnqYX
96tsWqTZ4tRMRAG6mDs0uQ==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
CNJnijKZjFkkzU8JHuPuGBTpITixwh9oXpGyvGPeqcnKWVld+328SBekmn/3VYKU
1d5CUV3pnhWSBzEBLat57rvUXDauRH0QxFul3C7qGuWMa+jhwJrGo5XdMdKmI7IY
POFmKI9SkuWqs9r5Tzdx7hmEQHmcT2wXi/b2oxbVRf0=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2592 )
`protect data_block
WKf1ReXikcHnWulDrRJarJF88Fcnok+evUILI5jlJJhzzK0Kc8QhGZW9g8KlSMQa
fSRis0f2O3E/SNoWFsBMSNFnS0Yr3z8bbJtyQ/XZm86BRrYmdjyEB6erCp4ZtcYr
xcG3iVaSNZ7AUN0aWZ4/hqYOOvQrFyrXcqV/YmuWtCGapHqbP3AZb7qd18yNOL/H
0TT2GSc3qM/Aq8RN40tIjMjoiCfyhEjLggJta4eU4FU2XjwpXSWVLc1Ndt1tVOjl
sjUZu71SmNNmJtBvA+hLEr/66m1EhjvXG/YIoEHTiTrCy5CF+xA26IOvGNSx8VMd
osofSF06/rOP4/Iq3PBxQV5T4xkVFgTT/Ye1EuMUuEBgSBS/I0Q3Ks8olmS3lai+
wthItfMwt/jKfbXj8Vcv7abOLiXVVjyrKuUMO1MJcx5Ho+HU26t8rWKhM6PRH4Em
yR3t7BAXd9G7kHe5xDB0isadk/JGbPEBEk4w4gRqXbAK3AlPZ/onZJ2bHPseSz5P
BDjmvUlfxoEsHkWy/Jfa1PDX2xbymSpk8OFxD04zNjjihSDnBEAOYZxoH6B0utx4
mUNSRhMGsTu8RrdSYwOuwhQLUihRy+HrnMiMLA9JREagX78Xq1aH6lzwqsVfkvDq
+K2R0sjDSY6DW8DUudGSTlNjB231qOcJZqwfJjUArtIVfS8+nCLRn48Innk0MO05
82k4pEQ1ZMiQM7I3k4zYgzy6R9fEA14fvQK2RlshZYQ2SHe7U0UJRWoK7QU+SVwt
hkQliYP+FndnWsp4uAvVFAn4XQGzoyG6ROKIGKbdCGCmOJTLP6VoY39MF4//IIa2
OImxTdB9kny9tQ1pkoB3ECUSZKvnJue+yzezopvL/VohHs12SUutPbfBFPr+6dTc
XfTfEaoViHy1Ug9m5Kt6FsHJ74eSd0qk5EJl4z9PWSu30JsgUNpp+Sp2rm7wx6Ef
fxGsVtG+CeqcZGL2lfypYu+Wbc3XXBV7afLmZRVMZOl2TAjX07f1D6uObYhXJke2
WJvbckrp/IO/HIVtWEf2icBMaccey8T7MIRwaYrh9RHvje/DkRofcUJIekQcgpe1
k96iqmHkvyPEqrRyn9b+HQep7bzRUaZ+oveACyL5aHLOLMERobEg6AyTXN89LynO
cXewZ3wXd7/wHrveZ/upTzsLMOgYOMklwrl6z2vsuiJHKrDNhrHgKTUtI3wNibtO
/upbjhhArQSTK0LSEKeTUdlsUaECBvmDwan6QTr2HNQJrNM9l9an+7sIR3bPa0M+
AzMHaBP3DvFhoUFlW35F33DcG0n3Q7EtHvd73Q5VXN6OSZAIFk+6qk7EPse/lY90
7czx3kw0FBB8s/KVwVkoiQhXl4HUKjMY5tn8ciRJ7wZhg5mrF3IcBmmGmIroFiiu
ZL18tlEXXsvAjEfupFtNDXJ645yMxkTdXhPoYzpY0UJ8jAnKYzJwUlb2o1BwXLy8
C+cT++RXDv/y4Iqp5d2jYsdXGHLZLPCy3StHfAL3VuKALnlmvZa1yDmaFXcDKA7I
ANM0IyVyeCpk1B/n7x5nw2+Lkgl/zqLdh92EYQPGxLlHIbh/n2lQ/XrXm9jTi9PA
N8pmppPY7bB4AXt8Rc3vNb4tr2GNlyzXOwi9yaF00W0JJbmpmbvFjbKYvNjd8BZD
2a3MMkdqUMe7pY8ua9ytPmtXn1ImI1IqIVXE6f/WU/z5hR3teNjDn6xigSvenQrJ
zlir6VUjvTX2GK6HNHV2k1O3gVVHi1U5CEiTV1YyFH9sVgUk3ThIjD6dfNUCPd1D
UayqYUVChSXpqpwzA4I7Zwy6eTyfwgTpWp2zd3EtHKlqcWUyIvKODrDuzhGrt4QH
uq5LzoxdBJsqrZr38NcpsPZk9KrwuhgFSSb6mZyfL7DbUblHSVXvg3njDtQQF53f
rPxmYyN30rpvPpCiIbokJWG3G28pIZQqVSzVyPPGvI7Nf7IuVVBahLzDZkyeQD0v
wU9roQBw38dGGe3JNxS7uMNIgLluI5mtULYtXEBzKYudcaCRN4sSvzWUsyydp5Ke
NCtbtBM/I+v4h3oYIoq+i7lZ4Orus3twhbvZOp1gQC5m+HX6rA5COxG43GAoN53T
ml2rcnd/MSk9aiuIRu0p/qEYk9SKM15vHesHHcT0p4nqHJBi0ufp3qeAiP3VxStr
t/8OXm//THnQlJLKkWPLlRZnBMdzmTDCvCpy28v1+UG/dCHv9kAojQ5keNPQ6fiW
tpfIk4dq4wrZMYlbUxRxK0uwJXEkN6y7o1+GVvZdsCKmIA6ZkxGAdc9Y6xzgN5T/
cypNQvuCH5RJpziovutT/wP9laV6Ndc+rS2yuQP6osiZXrqpMCr9c77uvajjR05T
nXZUQ6TJ52Cq1TpTZbVTQyJqKRcyjGoGyprLK/MtRK67wC2L5XP5cEVaHDIiN0RP
tzFAeVWdsGYZZC3Sw0mGQyKo2ZmKjlKt7RomQALhwbNP3S8jeca1Za1VEVHvGIrT
vKVCCrFWEjCeJlrl9j2l6VVqNJ5FAsbHaOQOVkQu77XA8kzGTFxjMwpo3EC1Ko0m
qLGCOd4CTfCCpFqkzNt92/NkgLhcOO0bHKxPCIR5qsqb9W1+Sz5ltTdjuThmkgF/
zZmb3WsSPNDGxxYyFPxh/6vmG4CPoceLfi5+V9GTWanuF/rzSbOJ71fhOxaJScVx
U9qJ2DcsHqCfZeCvUNPRgEBf9Yh95smgIXzCmOVeZWjoPPo+pf2OoNJTMra+Flpb
fkcs9xRvDwIb0BzdBc0MlUDMc+HB/IOHIB/4s6pKYFejSPwIxC52V6/ZXXBh2D+v
i6iywP/MEqZZ3BjzhFWqS8wUlEc9bHotWqaNvUAJ7tkcOb70h4iVv8KT7kwMaaNV
KePtGf6t7zojzQehtug1bYAc4fF8dD+R4n/W2HmtMj9X0jlRe/2YBgmW6dP3xkoB
j2VKssW/ewdseW7+5zxSd9kIu6nL4Gnhj3kkXSQFIH5zhkmVJfl7wuUOv24/gqpV
1U8N1A4hAAOmHzifmO4sKy560+5Y/DSKWmGPhdWPewl0nlZUWQHhwGKQzOp2amqO
nzPxh7gVe1AlRQBrw+sdOcIgeY3V9batNnUCU20u8DJyVCsrPttQZ/vXuDLFedjq
/xfFycR8ZFm5VbEAtzEHggBfbfyQEmunMLNeB3EBXC5mepcUra7Oz5XQe9+Ue297
qU3oozRbXVAwWzCpnVzzbpc+48Ps30MNJF17T6fNxMljdN0FLvGb/ZjvcJpibmD+
BaTXJQHRQpgsD0KhQr2hNS/+bwtYtjK7dQcN482w7D8IdDFcENArs5hBu/Ygu4qz
AMysa/Od+PzF4sFOtM3HRRbps4EmZ1Qkr8B4pkXzOxEyemwOwHSpfh/RjIeJ5oZM
ZbE4F8f01wMddSt7dcDFj7Ud0ZcHcYLRt4YrbjHSNNaUI2seM4os9nbJYqhnxERb
`protect end_protected
