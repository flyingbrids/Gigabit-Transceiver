`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
GAqGw908T06Z/dce1TwErCEPKq6Z+6cicMPkaQxvC6QyT0x6Ojkx8YCvU00MHd0R
9LOXE45IJzjSfB83oID9hm1KQB5HtwULyL5n1RRqNbmQ9eGg+GqXkW8cCNd1HfzU
jIQXlVFON2TJ7LMUstYN/OWJ1CstCYR/ILwHkCmg40PMiwm+HAH+h7C8FyL0bl8a
pZXBCW8lP0SN9W5o+nW5JunxN/FY4z0tKjVy+itVGJWOlswUau4kaqocvIgaIDZY
pf85w/5pplziFb1cBllApG+yqxeJcynluZujNhlXxZ7ujj95XIuANhSeThQEBNVE
nDkVvdAVlRXjB1uzcwC59g==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
XAl4POaKIVF3T5dGZ8ZiufqmzUPuWDdZR0uKcYt+4IG/JWdEAvaS/1mbEPW2aoI5
Om+bMGNGkrAgK89FHmi4Un/UPgnG695ypneqXoDo0OFpJ3yIGxJbF15f0/ncgIub
PuJtxNKPdTR7Tx0t4Q5iVVZ3EJoJWFlTxIEAmw9FkuU=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15168 )
`protect data_block
OM7pUg8L5lI0hFNXNW1oKZfXUofmtaNnMh/VSjjKsNhMRbJx7HtrJD70sWx3XLMw
W72VBMBhmwMGAtgYBNSpXfzI4TVfX4XtM1Olq+iNMnlHUt53DbmBotucfPyfPCyL
uhW/ChXm0mWHEkJzem/1DmRk5aWClHYbc7J7I565gJJOLfV9SmKY/WagMsFeOVrr
dJFHmmoJTi7rrQceAcNxZuTync4AHnsf9mcfMKoTT76dw6OdUv8Ym+7EJjnRF0hM
CpWmIfTkirdAskLf1egI7YyN6AGWXJhUloc+zDbI7YNJvjvP0xqiFJiZ4s9lEPYG
bsEnG7KXNTGevw4oXN8uc7t1KXmakEg2WdqabpDe2H5FjcNW+xWlfeKlzIhvpWTp
oUnsQD6CFNK/nfWe5l8Z8+F+oYpzc0h4AZejZRz4gmVuKMbuC2/5SYDsViYBN39b
v8+pfunO+HTIdeq9m9SWKVAvG4d9PHJ1YdCOrEL3qwofUnmzooo98f9WATVIKR11
EA7HeNPX0yIy+sx/Zw8tZSw8YjVKeh1FB7LW0+Yg2UmJ/EeA/7kS8piEGHngH0Sb
Ne/TgyZ5JaSEoHcGYFM4KZlL9/oJj4xQnLzOU92ASZiAmmoVxSDgh8QTyvfZd0F/
xUmoQbQpDY6ppsGXzLUdWRUst/jPQ3S6C2QrE44uhojfUf9yl0UPIDP6jPCLs4m8
euP20dMuK0eNW5a9f9j6PJQou44VM7YSvpj5eC3TUTfvIKZtw3niwCvja7zjM1tE
GgJY6Ipf6Wt8czbxaDVNjkP1Ylx99PcjxOF9Bl2jmHacgVzR4LlW3EvZXZa+GYRv
b9jfUzmpp4oe9eH+LWRun+/dNnCbddIMygWgx9PESvFUKFMOT2Iz5AeyVFRRODgM
ZhIxr9iursQie9rwOlH1unouoL3MI44+39pk8F//0j081Af0EyfABoI6d7aZPe3G
9I2qIYVd0ikdTiJycJjTjiNvNfoTFgDZPlutDQxizvIgYgbssHBCxrNjkB+Qaw5k
UWfsPBqmeT/qqyV2OXjRNZQkX/AyEUjnKI1YusyRojzEMkK07dqJuO2ORivOTVWl
v2de8lLHJ4ESC7oF+j1sBKWTVydxEvjsLup2BeQQ0UNcjHNHf5KJxaAs+IG7luIF
HxK2seV8IkOd9qP2mNVrBR/ccia8esWx8Prwret7alDS92MFnWP/AScvDaLGLQN9
OdEffC7hIy8exVfZNNHM72EMMsmeSAdO9dIAl9algT974XsGDS97/Ic7/upsUPCf
gxjpExMqyTuSCuOPXkXsKxstgSTPM6M+d0sM0c8VGWENM8TJCpW7izAOHFXJfDG4
0hy67eLDBUV5nsFLSarOc/d6Ll2RjI5dECxGKnmBCnAGRjGokn5xulLzoPwV6AIo
2/v89Aagg8iwheN9rcWOkoNgDKbYySEOc8iB+BKUWlL1dWjd0Tflej1snLPeoNwj
EWS1WYuBgJsHaLP60We8sEVxCDhuQDBy3feEy67/7TeNncAKPnsHHF0WrX4X7kLO
MtBKa8F185u9M3NdrloHK/R20rNScsKgJ2oRW8SepplyCOZgJbf1PvjEglTZWHe7
unSAJUpZNdiCN0JhfPpGgWgktmfzmgzzw9n7SZBHBTta/XxCdjrlkrTqSEnkQ9Co
dgMmm5XQzjmYHNeadwNXEXSgxLbS12+4qJrZmUejDjPuZwps97WmVvY6bGKcKmYu
jZxk1CS/PMD+bXTQz4yjzxSAPTI4uROCO/0+0ibOLdo1NV6ojWJ3zHtJEZCP3tlu
bdqbksRvLJAQoBsxdT5DWonf4VmTkgffjfX6eAjrNGuTLXmpCBV37Msy5mg9wzIw
C+jWYtvi2v5TXFknxNQ3y4iUAYQXeXe4CHEk6pRg7paOc2LkLlnVq6dWAPraRmIH
G/lEAfIIgn2JUr0+TAGD+3gjG183UnzI7uQqZ7ZHSYPI9tLipDUjwH1k2cHWTivk
xFUQnT6rLLmlU4tnTTGAFFHr3x7OYsy5ElCbKAeJquJBotwVfSDZTDtg8PyUVHm/
nrM0UBznAQggKYJOZJxcZcnUXUmHbGIEeq/0jMN5HncxnmKbVqnpkgD3c3ivLg3g
uY/9dJekPC758PA3qZY9YIXYJVeYDYCg01jWz6jBzHFHkmNL3w5eXP00pvm641H7
fMLvuBqdal4edtz9PUmgYmTN/2wgFkFY3Vj9jEWYGfWrYR62iDXbXZyHsbuXBSNY
+L754XHGf2cpYAem9G30+yknPQWmOf4HZJOIbL3fsN8HdmuYEbHWo9oq2RFCr6p8
NF6SEVhITS02RSCwKcQVeMAexKV3AKaq356ahci4yRDxdO+0Q119Jd1pqva7l9aO
Kamk6pE+UKuV7009RXNAjUIdL2OeEvi4aU7eJZDGPxbMg+p9BUymYmg+TgJYmOZi
RPIhJHT1YAypcEfdw1385Lv4cShvCPXrAe2VEymQT5Q3ckPg0LX2cffizX8cuK2o
ZnjHdiQ2lMo9OIn2PYQfk7piX4vbmVygE2ew1YKpDijAQa/nL79Zl+K6+eXmb5qc
4c3EFXptsRB+yUfwGMRmVd8C5slCef+JMxCDtsIu8aQOVlsNiq4hFVAWuQPi5zV4
k/3Nz81oVu2+U9/q6buhFEJSegQjSpBFYVgvM8deG3zRjwoTzcypdxHdnEaEidE/
3H7mMZUPDOExvT3+GOBn2fO+7lfSQ721oQ68Z7v9OJCnUxIZLD8lKvLgxQ3oyJVj
kyepIJDoT1t7nz9FZFTX0nsxjSj14CV9avk0OG22oKRVAuy+Dq4eBu3AwBxDJ+Le
nbMAXPxNUcSMkOyixaLVscd61p++W8NlNT7yqJ9DxrlI8B67k3AHOecIyRDQJ8++
BF0uqFCdNWQ6pVSRQHXzf5H0wz6O2fikw3polCj6YPfulkKMM97LVHuW3AMLuP02
aGYZuIM8i79GuzRDZ8i69vjpD+SGZcmRrNFalHkzw7Kwr7JxyqUR9CQGdcDFjJKo
D7LaKFYIY92JtB5w1go5NpPhNIiLt7tuW7qqHLnt0ryl+HvluVRC1FYcjf+Fd8rA
+AXj6gpDR2o0QmoFnSbA/SDWLNoe1mzE9MFlWXzOaTEhh1S1yNh5tS1johfWX2UD
qmym3ScqIAV0zUhGq9bGKFCALTATBHDQVVGWCXMTZlPpKVbjoRh0E1MqN+FP/WG0
0qII2eDIz24Rfg7NbXAWPknyMtQbDUfu5Y18qmMl+fGNb2Iyn8Bitwap/JwKNlmL
u2d9x1IqxsZlcRDB1uuiS8ME/d1lzG5tIXqJsmJbfViS93amjux91Ovzha4g8MIa
u8Z9X3uiXjq10mtX4HTYo3wXV+UHM9B6cXam83wnKiqzPtQ+FM6R8/hmk4wdNTiT
UdXB0oF4qTBAdCwLQnPqpK3VKc7Fvmzjjf4R6qqc+DPk1SsPd8VIC3qesDnZQXVZ
T6VMnEK3PEnuNcgzyW/FyUm7XFoBINwIT0VCD/nm7GUaK9pt/FObPUTt3l0/tuwo
wZsooXI4bh7jHaJHShb8Bw3C0M1i+z1Gztpg4gzChoiU68zwxkU472wzIGG2AX7P
wr2fKIY4xKDN3NGzlIEHIJvA2EtD79jIueMrhLK+Cg7RRwiESv3vx03RerCxIJ7z
Q/f6m/9oQ/j+cbthJ5OdPDjveWLGu6bemhtHum2+2nrNQuQOWGeEDC/XAIK3MA1U
pRlZ2uqCyO/aOzygrVyPDz/CWg3KduX6I6mTHlFw0cUSnfSzosEcGAGKtfqY3rZ+
k1EjcWcsIhnCAcnn3z6+OIpgOWY7yIpfdWp1FVBBv5zWR/9h8BNTVGeXj8jzlxDn
PqE0N+NLq9MkeZWjMwvx7uCvQ3RkHcXfVovWH0ZxxhiegELGZIyvvZJXMNODYLhh
H/NG8bdRFl/OSN3vIuBq7BnAIuXJtjSjRoPXY2tRpmYKrBmeOJhatj8KaBztFy/Y
PI/ZzkxCiElZGPTFfgTJyzX0Z77dzCeNB6qS5/7EzpzufodSq6gStsdyjlVhxNZW
bH8drIX+NPzJ20hBvQwTU8A/ila+iqe4Q81BbLUwHNvnsT2mVuqBA+uonpQ6N59T
LjM0X9XR1rnAbv80RWVPpjk/YiTfS903gfMhGZVcC1v73OWr7Ce2sLuau3i3dltl
K0iI1fzZzgXVU0cyj4Zlb7S/VV87phTCqB8/NWK0T6d/H+PqkFyV9f2eyyfUDMc1
sJUARFAEjoprl2hsvm7jscRNUY3nbaaj7Wa+jMqVZ+9huqJ+pVljQgmQsdGKwpEQ
3tnBuJJkq35YAi9IH2NUXCsbOa0mjRUH/ZEGwW1WrA0iZ2ucakiyjax/Fp2K0C2q
6oanj7yY7KBAQFsB8cFRnwSZqhEEd9+hs0Kv0j0PCeekLWFVGcqu7V/nflCwrbd+
FF243cmKtSgL0+Ue+uBZfkuY1ul7CjxMwvRZ9kd9CBY0m1XkCI7w71zRjthpr2pH
aQtkz1i1ID/J8zsUriPbRci9Cx3KtngHiXGogGnI9lG4FFCkVg7paoScLWnjrkZi
G99SyOfBO5XWjqMVepL2TnkkeCmLqk5tfO7lIg9BluT+ftWUX/DS0I7wMNmZtjV4
8vlIwCknlNyL5qOyshOjh+G6oUpd7lFrutMpyKLj8PTL30DmU6zMrOOyKszdSaYP
Q/vK1K/CVexboB5Q4BTnvNT/MmPA/38a3iX4QsXfIMXdRgFs9ZZIoybz05Fg2jgq
JmiKfobsqwr2q2eFkuuPtI9M+o4ag0x4G5+gpPbrlQHvTwjjmeZ31+hzTOY4jYFx
Y58a8YQxPixCtNxIX2aTp0H7hsoxuCmyCf+1gKhKcjrUYW/skgDVnjH00xdmhbEr
K8sPZG9NvgvgMK7YzaWItF1BSw3zWb2Xj7vWa5Og6A11I/TLmeaXaAk4TqmfCeRc
C2NPh9sOPa8GkNpzPIj+7bFlElIGc6lXOR9PvY4QHVbswi2KNeF5tRSB6A/7iW26
ewkV+Pb29INcFyJXykYfjG9ZJR7SoNKHjcf7I7Z1aZG5h3jYCCoYc8GVVQU7Ccoz
0dRUSZtO0gpCRsAVOrNP5o4KI8mPLhnjvoJPKEN4AcsS+SlpQw8itbaWRpcinuyV
1Oou+GFY85tBDzlPAiRtY80lexaLxoILNipw9k+HmEB/0yOFQ4ZYXXRHii3ks8ok
Tvqy1RaCpf2hfIW5pRDxpzhCLrZ7xoGdniSIbaurumbtkbU+LMeTmuBIsmabvjGG
YnNMtu6a/hmGsxKMyLJdgkyKrDqAB1CHrLAgUXYCQdAduGvbdo5ihBc7Se0pRaDU
r9/shmNbtbse1NfRrozOG77/f0AEuofBn88v2+802FKxV+ltiCEA6sfJVBUxZiWf
+hhpSeD3cTJL6TySM6b4/jSgyrLLUcmrxGFSi7z4EBWAIfqnBx3bJZyXrL9r/+pq
HK07F/Qm97oKAD1y95EIUl5fvdLAEexw4wSili+PP00kKKLGOhcczNHlIZwzuu2N
aj7Zwoiac8xrDw+iEgATaBbYHRK6Iw0oebqYstR8FSF6XdhBiLM3X259T3iG+DqP
CTHGp0K70cDz3ddlUJv7eLi+/SYTVVelurqdDXLCRpRzBzMNga5gEimik/9fdOkA
i9lMcAjjjL1uy4TGoggRPGZb/f/S9iMkQRXQ7VrY/8tbqPh6Lo7X77Hs0PmKyOVQ
UoeisBWMZ6XTP7i5U+17T4WbRNHRvMN2ttZgf0x8Q+xalWwgmqRUR5GqZh/dcVPv
IMXZakZTakfSmN5WvdrCkMizi6YvPOZxinuiUTeVLbP1v5zKr+u8K7scX4gPoO6+
22X/csC33dapJrEAPrck+wxh3sJeJFHB2qgcr9yClKvcJhEcx+J7diJVPZxbvltt
Q8nwULfgEPdqCr6qrb9WPVskifCBI1XtJkEz8T6tMzhtOqIqvNrcCMzjC3I31qdx
9hd48qzqHlfHmF1ryXoSQxSmDyHOpA1L11fiF4pu3M0jXEZCyz8Vy0RREIKVFns2
n8pWdzBVXDqMsrSZmC+wvGCzzIrdTUo5C3R1R8jS71l/O4PgG+wUjNJzmnC/1eW2
Rk9TxqcnPzJF2oaV1cdAhp/8v0ov1V5DtJC87TUfQBgL+Sj4SUbuVgRSX5Zk451A
E73RN0pjXbAwzPtyl3MfUMmzj2RH2PvENdLJhdTB2UWpIvvK3pXzXQ5OW9IIWmMj
dRkeiKBRsH9zITL18UPHx0jGWlGOtsssp/wjDrMjmbF5uLZ5fmGiRmX2kzF/P3Ud
auM4dwyQbo8fUiXAOyK7+OvCQFi8LJYGGkje5NK9M0vmKX2qsp3cGuHIcZ+OHt45
ADdBZpYftTshtb3dgloRmQRiA/OXs7n/UDJo4q7Vn826wNipDbppEhzqE8fcZNdg
MF63D52t18FWX9A2eFgMKQCFnoCuH1yca4OoeQVP789TnbpnIbnmWJfZ3o8qZe+u
xQAuTNrz2xgu4AA8Pr4aWj3s/5KYFWxGPmYyx5TTt35A4t4dza/OBJU/toJy4Edd
6mnQsVqQBlpxAMRIbTSYNNYQyKJVzyAzXP0WL1OVYZiDxnsk12PThouQ/XwzCLpg
yzWmQdYOgjeCOreIZ/eFyd2P+wymlN/5iQUfn6kjhEq3Vpk1TfFmXAZxC9WZX5Lk
Vrv87DMXLtUycbw5RZtreV5a2CKUsK82QOFfMpYm8S7JTW/xLt8yEQf/x+pLxT/8
FZz32bboyHY4VExEes0D88eH0wQmoB68HZHdAp3oQjCCwevdeGCZzxNzbkqFjbW7
ndf3RrXNqDKfRLCxWaY+av1h+76XDBMWLfmpg8u4XUjPJUrYK6VZFHJ5m3K7Z/EN
Y6sr8JcVPLl7BYIIQxpN767ccKooDcXLmsVUdER4e/MnNWL4FcThvuifBz/Z+vGl
K00gcVZmaTU3U/a3NWo6Uwg77LF8AB3dr0x+YjrRoIJyPmV4rgxOOCfzo8u6C+Ca
lsEXcBZ2CneTJmhIc2Fkp4Eg0geZATXiAS1g80cuDrj94fDYAkppzoED9zyfX2Uh
UNQ/aXIwLBfj6BtaVIf4jrn4DkJkDnhlpG43oC8voUqaOSEtnFqwHlhs9bFZVzUE
7PSBwkZ1I9RZnimEnnIvFOCZtRARdlxhxdxQmKtAhFWJlXGa8azAQvk1rFDakZSn
8oSMA2jCvk/I5DtmIiUAzmSJGzQ7AdMeGcCJkzxXR7i5AX5I+MbjTX9YQ7luN6Fm
eK3jM7ZSMD2jX4hgXs3zUPZMTSmqcdtykRwTzqMYfqk8DA41iw7PxoeujY7DwhAW
1ULj5EO4k5ELvGVytdK7duu0dlsWiwXIJzCYXbVDFw7+8m3/UZsIFSzbYNhLqFVP
kO0lJaAXYgfGkp8uxSxmvNalUBfLvN7H0T0UO+qHg4dCktMakSx1aX7CRs2bpPMg
2yQlfE+aDZnT3sNO3IfxwY8ale5Xh4xMWpNXZ7bXToyfHCy28wJRqzUAZHCDMLs+
eRz/0xmlKN+l+X7bW/Dl/kSUULs21+F7NXVg0vpF9i+MP+1SmUWapwawKBIv/QDl
fTJb8yzGpkQZVPQZlFIjv11vuFD44KllocdfdKoN/8oU0LTfRDBWKTLv48xj9iQt
FWcbnqmyfyc68TFDbaYzzpG/7YLW5DeMEULQZAgJXcadLwZRPkmOHgnw06EPdnBc
fW7/uzCU87eOCSctfVx86cPrABwPJrKpaiXz5QE4OzvTkLySIwoaP80YTuL0/Cfk
L1Y9BlCp7CrR6o3y3PfO2eUWBNDP1GKA91pk5jbzGF56FwEFqItNqjbt9juLvuYs
YJeI3qQsq+G5rX+Sdj3KJbWvz5qvirtEsN6lvWLYMTLAq+dMjcVAywm7wIX8AVV4
6/QkJWTSFPdlMd/nj5joMSg/v0aOVPNCKU9mwfi6eaBWUFJaLF5o34QPBRSqW4EW
dnjgtNyeL6uFlfng0qJuUuMH+W9wHiOE3RB4SsbsEWrFJkhQUa5vvYem0QWAeolR
PDg+z3nKJDqT4Y1vY2g4iRf/jTEK8K9SKRi9gHCK0d5fx+yD3I0xrBPFhce2gaxA
tWGz7nBkyKuOHG4mCNLIi+VN9MM70brviQ8Kplov8BGAmtcWV1wTZheqBieDSbKl
cR8VNJT/lmMw29mxlhxl+bhI/cvcG43dFbUqtJNe6v4bANKU+1eTT8P7BXUeNvvk
Sv1Ki612ks1CxTfbEuNXNN0bySigxxwgyn9/fTAKhUlDNAfUhN/sxSnkEU/US/vN
m9HmuDYT/EZkUEE5GgwEBSsMt6tjV8uPO1ucfmZL0pU+ikPs09yBghoee+ioN3gp
HAjS/ETGRUNh3gG2VG7j0hci8r9cLQIu7xoU36oBbN1ml/YKxrizXkbfj0KRqZ+S
SkjTKBgDXiC0ZDYLIZfX0jZBTxYpL7D6G/PRmYUQfPDmLCjBdT2Oeb2FzYa2kGzZ
bCWjpkSqdTF2zU+1UvncGmHcRgIpWOAk7v2qj2UGed+KbnqSZCzdUDFrgFrIb4pT
9gq7F6+4+t+2wx0JeryBuC77NpjjNBLQrFf3z7pR+8/YBisnz0wyjhkdPcLKHO6R
gUn9BHeIGlXQXs3hqexhOk8y7lDLiGabbHKkcGxIe3kAWSsmqoe7xDt4UmsJhz6T
L3wzEuDkwc6VWoZDnwMQ11avvo9twvifemHneg9RhEbjNbVHdCaY9LR6qqHeRz3E
XKh6aqvEBm+7vtqVPSOs2QSxzxt79T3mX4Ft2eufhF6Imp8X9+XWC+G9xpnHdGEh
KtEOPkoajCGO3zThlvhGEThZhyMlH3wAQOZ/gNYhGlhS8ePkSwF4vq3zY3jbiRY4
dVOi3LcdMOisj5kZPauHRkCyajB58ddu3D+t4+b2CvVXxBUi1f8V52J+KNBT0V0Y
4B4Mcbx2E1A2vn8rXmHHfV3cULFVtfWiFsfSEf6B8uwTAiwGC9rZ8sE1cY5GqB5T
A0He8kqty+edNnbVnT+x5NoC/Ne52xse2mlIDUGvPN1sD+0YlvEDJOljNuMBr6iN
EkvBLfX1ZqgKwSqq7hBdfIB6vHvKOfAuDwYws8zSXA+sK1vNUwaPmaByfYCKF1w1
PfVIm1GdV2QFqhxNa8NYIOxQlsjWW3jcv4IDhsg+8FJvlGlcAb7hdQlinClZChkW
nGdnim3AIkbA2JXpBYdW8hPNrQ8dawiaW7j5/2BQxCp2DXL2Ndi6KMMbpG1Yyatp
XF85uhBo66wSbKycqahbL8NwuBxqgRYyt4TFFQPKBG595nTH1ObKqMLg9Tz0V3N3
op/wq+ybG8QQTpcGyu2mNpWwdsAemEub7Lk8cTIiV1ZsTmRK/K4dgcS1d3oqnC3N
MHTfOVAEW1IYstz4mRrFS780ORQsk46VXW3EGhnpuyNZPi/lY8eAGTx27uMLBXtY
pCth3p9FHvPYgA7nnCB5/9scBWrEQ4wAHnjK4KOIL1PpBUEqhTxgd5d112KPD7Pu
1bsbsPl5q8zc5xfyY1U8AtynS1EhfJb5AQcdcoqRXwDkgztJHxPi4xmbsrumaAZV
wGa2/2cg3aY0znbPiQNbcRtWOFAX5Szv+YXIIgJ2WxKjki0t7LN3CHfT9BM97bHI
pqdShqJPfeRCId2A+slVQGLNzgYSJ6vPFFIw1ODJU9ZrYtmJZcd8kt/5rTDcmzQj
zu3Zq4PQABQyQnjglgRLYsEPbD2pczF3Rnc/3Rbfv+fVjEp7Z9+6dLlcYB1+b8O/
ZhnEtYGdJ5vQYIy1g8Fkj7n/Fwq4WdGlpl0C8kkBn3smDnK9ac6iTXAKp6q8NkmJ
s2hCPhPLDihCNK/hv+EKD645b6Hh0thviZ1ca7JrQUWrsNAQOOBe4aizHhs7uONz
ZpVgEsBmM3ciBQ0YESHwbO1P3Nds+AX328c8Qv33WcrOEhFTDddiXngUE4A7mgCH
2sTLZhqT351asvcYUelJJ04iunIkXdqQWlz9EIBmomTPxgnl30hdxUZu+PYgphoy
To0TFR8qi68jGjLZhXPc40PFXjYVCN4lvp9BIaItmdFSkWMVD4VvUcjiBhSUTuLA
SetNp9BympfvlVdBFHk+6Pd5Q59GG0bu3clVKMIwyhGNZyawoGj/eL0G+BGzXIy+
b9wSPS8R9p1GGpbiYK2oyXb3UZZCihuwLofxfin+pWYqybk4mXUlBZAQqdVMeINI
xFDM5L4I2w7mMcwnadG/YGNy3t80/s/p5HxzZ6hTYJDSViAlmP7fCsoXwYLg8TOn
tL0FSKOmRetIPpS7ISi9XpjE6qjZzGpsEcTFhH+OH7+Xb8NetiNb2dhRibtyeo1p
8owjDmChGT4BWeoN9zyjzDDCEyFgsSFldjl12kRRzGbtKQVQKPPxwDRNCfy0ODHU
WHYH4L3mB/SK7WkXXavDSBj7FnXknfPxKDYaKruRbH8LtLZEw6cvtptRyWhpVmt8
snpRJ+Mp0WQtDTEKW8sfIzRvNLBuDXXa3gL9zpv6r5rYBXyHhOPQVItHZD3ldOYb
D4y4YttV+DXccoNHK2Flfs0otLY4UQIYZ3ZFhub39kVqcx9JixP3RlomB2PH1AmB
ihgou4YL2oQeqxxcyqYjTqAsv7/3IcDR3YJjjK7JNDBQMNufONoLSyV/BzD/HXtS
yHxOg3s+FuAx2Udq9xCEc4K1xzAfxcKzXLgzmLhkUyUNUIUPk3UcdAemUNeZ/dls
JOuyWKkV4AYtA2cjLZiCcLJPHqem3vBki+wPqqgl6QSSo9NQbZZVvkYYJI6CV0mI
iK0qcJ4JxVAf+bTRouSYOY/vzlHenAnH+S47Q2KIhxSC72edv6aO5lF7n9N/y3db
xTTvsBPRm7TWSpSig2nkyTa+J/DvguwA7wxlFoa/XKrteBhdl+n+wy6IrKw4SVhx
W2hhXa5zxANFceoUp2PS7bEGqmj0uOyAuiaSop8IqFmJ4leH4uLyHurJZ9mmhYnj
2FuGwZcnxqvsoZQstlweIsgG1UYMMOImdL9pNUqAtdnjQ7twpQIpwoGlAYmuhN3J
Q1t3Ny9xRnDvQ/UyRU/u3kwYd8lFV/9LTZW9I75QUmkYB2yLkMNS98p4flbzaL/M
86fKgQztikke1sWgEq2SUQ3iftSJxyZfJ9DijUtb/R6fotwOwWk7ff88BoISeSGX
r/arnf1UI1oaiJY7ELDmgCJVTq0wChlHiRGzuSWAyN+xv5p1LAOfagAsC6/8V+/V
LDJzBhUbLBwftOMh7iOOSa1ql6GBFqS2deWYLDuvrqXu59QvXw/t9JhtfT7iu3aT
GqjYH4tELD2nH1LUFwq+2gH9HJPzUdREtaIFL0U+NKHDsHQOMN5UK5zObbID7r7d
7DQVa173xj6hMM/ghe88qcR36tp1j44S0V9ngDxQ750hd3yioK7QuqtBTdNFw6Jk
jqXBs65UI3aWvtlvfRT+fhsKQRbQDeixTEh1CEsEmhjyewYtsK8KxEajgfwUggPT
62Qhu7WoySfS144SeLq8Qqafs3i+HBy9uenxKJaB3Y71rqHLk/VdS/WjfoYMLrJA
XC8CVcZ/rzJAOHXMCZOk1pHz7nSUyKnDEnrQeyIVv9ECnpo/JCnmWI8pYa0OL/G2
o+wLcj8mLDrUBkr3Wf01sTkv89VG7xMmkNn3XR3Qul6i/nqmIPhP7ygRxZ3lzq4F
l9gRqLf1r+Wr5fzkm1NxQ0Q/XWbSyslKDbgdxNfbHIIvXyMUQt9cWHLYNZtG+6iO
hKVfATw8h9I0ArJOp/Pez6mG9aom2kivCzbsdyWjqxBLvjJZbFch0P1aflTLcINn
FttmHn8A9BCN2k1UQ3FwBhpMZo0a6nKrB4AFitw/TOQ6M/NsuXJcoW8ryMQXWkKs
VRJnDYMQyNMVpzxFNZFJXnH5HvD7oswvxTmEwhh2IpVw1aTjr5HZqk5FRhC+DoQL
sfD0cUyXYHNLn34W0XmKsd1U8oe83Y1ryistkNJEdD99yckFi1SMY3OVQyOaEBkP
EREzGWEBe5beD0qdrmCthApapsv7j+67bAgNUp26v0xnhFEPsgwOTj6hkUa7A/7O
kr635L9UWYvDmKpHo5AqKXOYthUcTNkz+gPCxaO3irTFI5ijy92tMtiAwhD2TEAV
YS+MqW2+IiUb5+EWZf4jAl1jU9TTVz5DzfZWCunJbv9ivi9wWk+jrpZohiSWdZuf
NwyOIw/6gym+HB9DSPlFrfChc2gyhoQo0wKifE0tTitZG93gU8IY1qPuHbXGAhhi
eZ0ugMiuifYXOBEH6eFkbRDDeLs3ArYTOaterxAjlGASnW0LjKXNfr79wu1g12m1
+4Vmbb8EfoVBoLdyzla9mFkregzshXbVBb0xf97noA67xZvhSM8aUhrf6AWlNaN9
0psKnEhwmkp2cGYANFgAw5i8rwGGEAVpnBOWEhkfbiF94llhRQXA1MumIbDAFPnb
sx/2urlRBwRvQ487dftkfw5eIvolOcbff+WvL9UQuID5XsmMFenjDy3JNtLKuITq
L97u5AQV4ggoJTh1Qe3tvUwnDkI0bzZwwGa07zBTSI6N6kH43zGn7OR03tPOh4oq
A6tZ4YfVZr+JAMWUV9aFJIfxKLuwbSc5bXc5RSPaphP2h+JZkE/hijtnP5pusRZz
dtciyi/yVZl1brhfUc6L/udgJqxL4/o/QCzV2rF+rAyuXElaK2WSVgqmTX5wG41J
xx5aljNiTXZYs6e4KnAzfMu1kttpTEwS5L3fdf6zfYaAbK8w8MJMy6ZlNfPEwFTz
EBDyt1/zRB7Ji30M0njIbORmvSD0x6EjKwf42JMxSQrqV3tAeEzFa4rAuryfoAzB
1GdChUUU4yzAMDzSQx23d/CSnMFYhuOkC5rMwS2+S8kmpxYRdE0kERcOK/jAf3sn
gT+XH7krnfzQsCZ16mm4tDbrx2/IQOPwqU//7ZYgsjuajb1ohBMXJz8hIu/4K/lE
e6/S7SQJKhp13Xx1nhge8jKotr9sO9Co0zG+6ljVPrri6Z6Iu01iBRKH/jzO8nnK
1BCsG3EyRxs2qaFDhjubPtaucvUY5a1XuG7E5kMyaWtziZ8b/TX/RrrqRUrHG+5C
Dttbbk18/SB9eWGBMw9phQp+cKH4eqFXOHFX7iqy6ZeGPwjkkjZMlaWYjfUYjQ48
/0MDy8fTndQNIBmEGY36+3qEp5kmYnYrb/Z7fcq+lXUoOyXK3BJVefvwB3JXPc0q
YqdkSPzBEQS1WJ8hZowsE3ghzvumupec53Q3hga87OHTJO47/HmgzgZImuPKRrhF
sDX1fM1bVE0gzVKiSxrrqU6Xy7odY9Tl2z8RxJ0JLThJ8tpom+vx3s9lKSAeRyoW
FRTazvsDhIsi8HThFcQvk9pSO/EfS8FD+9lTvatKE53PZMJ0C2MJAcW46srmGl9q
D8WDsGbunEv8Y0DpdkX7cVxAaV6uKRaNzUi1HyKtmnkyFMMuEmty1lvIfsD2c5bd
3i7ytkfG3Z60SlEnnUlgtju+QeXrtm6Dk+/WMdg6ywnRMPDLdnsncE2lcP7K2dxd
RT7sFBNNw77QC3Z0UucdA8x1d2wMllHecZ/oafdyXaWAl0ao6+X7x8owHfTbfMMm
Us6694CegpJFeUfxdXzDAhtFgbYu+gKNNcKvGUm64WP0cMavPW5grQyptAh/tB++
4HpXwqiLwf9J4Ac9uZy/Lwcl2YIisLIYhklS5S7jVgYA6FdDNi7MlWBVei+Zc7/I
ojPBUEnMSeJLo2pYeSG2j6Wzt8kzBZJg6Dg81w1m6UWwR65f1lMJ4/OAQ4Lfxk40
Xh2FB5Jguas/AAHdNhbMsEPfV7onStd8M/S/M2nW5d69mpNwqDigpYYBatcHn5jm
BjF9JUnDulJeV2aVJ32Y8SspX5nN6AU/H4Gns01PaDA/LX5NuLdfG9M0rNVmdmjo
O6eZEqPHSnnp9j5uWPfQ0OhTaTlfU9a3Z8l4uVhHZt0X7nv88yB/bxCXJ2LP6Uxw
fKFRABbsM95wn9KOw7tFfpzmRqc+DiWL9LSX7yQiqJjG61DETW3Tnsceottq/Me2
gWnTCaZkJa1gpCJvXx75jeCW5sFXDodWqm88fOVmF83m5MMtlASxc4dlBRFWBWtc
i48Oikr0kWrCe+WbLUTMFVKM68IVQxO62c4rZBZBvgE4RQWW1z1kgmjQqnaS/B5O
DA/C0TLzgled8s7O1X8orIn24QHqHG5xWC4OAE7pVr4rULAMH1gQo9pMZlm5KegI
YyytuBobd/6XANRYzsWSWGqxtqEAZGM0L1hO/q6R7Efy0kuKC7WOhiPDrvlTgfhK
noCRoEhDgVjbIGlIgu+eSEXeU4u6FQDzJVYsqAhlgJiJOlWAAEbdZpVPqi6le6qB
GMt1jeTHosi5kjjawLP98PjT52ZdTsDrQHDfuLQD2RQp7qdrXd+MsMZQtqRs9bAO
SjoWlBPy2evjCYViMo6fA/kxQKEpsV7/B9xafheAWr2AY9K4O+0XG8hYm/R1A2MH
0t2MiKPxylWpYntN4l1GR93uGd6+9wUt4F5Xo5vAyoUpJAFABO2zq+af6QPeCkzk
LmRA0d7zKDsvY9gmcIfYiPqxQbH5fP5xqIMsJJMjKxnKMo1zmE4uMHv0gRtBy17Y
5zzizTr0l1YtGS99/vMB0mhpgr/Vr4Qoxz2dBz94zyEwJq9MIDrTHgPqDqpToEbf
4q0YnquDTheMQOVw67KYgxiMeZg/yAQ/065YXbj1/JU1T4WhdwsPq7FgP1ZegYV3
lcFKeoBDggMRZ4CJzAGAShxO38mrHvLx0T8k4LEg7t+znm9wM7ZrkqenAvTZvDHv
bUFGrD3Y2eGXKAElM6rgXbGco9+tNXRsbC7UPodTGk7Zb7ZLHBZemTpzsdKbF7kC
QvwZO935NWhS9nF7uK5RH8SqGibcAX/tCJF6IXCEU2lUEKVd5ubApwPsI+butRm3
spuz8fV8STNqWqJ2eGPKVJzyZ3Nry0iBgkJezv3p4N2uTPMMxF999fIqOuA7iSm/
60lSr4yKhZzGF9YTpPk+a/ZENWDBFtuPJzup+awESDP3eEag3/X1iwwEmKi6BzhS
xiQjYBgqVcX8uPE6lf8Upa4Cq4qKSJnvZ+SNNhR04TnFbNclEpPwraaIjKO9e+Oi
lyHlug/M49F0KS4fmvu6vRHED5F6rRNgi0iw3Ec7tFzVAFiHyxRLUkK85nms3Fq4
M0+Q9pRUysO+Z+pPS5uy4ay0ozC4Ok1M/y2VZU/juv8llWetf6JCLrTi19/kEsgL
I5r/suspxcRDLn/FlnQBmnDAwtPWzfz++7mWgNhLlxGDr5lj8/SH+72S7gCcdkUc
Vw7Hi9QR8zg2uv0/yWDOFf8/OCg5sldyTH78nBfq356o/9ysBdOWaTzsmsI/Aozx
XNGGDtJ4QEl7iT9oIASIIZTJxAT8/a4plNqYnuSMZ/vLxgGDzDvtvomlz9l4mrTU
kP+6A8fcvqBOfJSv3b700OyTTOaaMqmtvPoaXyInOIKUQw1PrS/alxI5+ZFS9I2z
SWgW5Wtb5Xd++DMqHjpnosEIoqcgGl8uH1HRUzKXSP06GXxle46V7FTE/dSjk2Uv
TE7HU06g+CpD2BZvK5Zw6Y2Tczgs/hsO/q3/W/5zfANaLAox2ItZlBdJDI8ZGrO4
dFIbDnnjGaiDtaUatlGMpWNtr8qt+CZx7DHGo71BcSx8Tj8znDilj7D65HgDo8Kr
q56qN2HgtEtb1vaQ354HfzTOMzcAWpe5xWfFgo0vrBY9rU8DiqQN5VMFsREcaWdl
t/qZw9bhgbFFRUH1groBkZ0JMPZ5UkqqX7CGUKVtH1NLrPcQMxKJS+0lw7xYCZS+
6+x0VQDB+re0UUP6BYi5oCzruDMqzS9+N/URLlP/j29W/p3ByLNCV9Rjn0acgFzX
Y4uM8mvBezBE4FkiWiFgQkPc4D8ZMIpWiC13jP1eZOhQ031UUweOmBG1csjwz1Mm
9PuYzWtNusOUDPlVfQlxn0pGCCqmLOZl+svRJusAId0WwbobPssxmcBPvufQJqC1
Vfa/FgLmARAVxcMeoM29VGsBeiR+QIBZpUy1XgBkbloWb7FhyxqXLE/cETkgKsgP
ntqE1P75vULQy6Wv21urk1c/5824Dw6x/EpfuqEbsOfNDvvRT/ZMdDRnDhNKLkCw
yZFsrOAOd0yD7Frr3aJ7Q1xuxN12BUjSXXinUeueJICpJe/2DQoRflkdnhHSVFrP
k6j0JyTDkRbw9Mt+cu7zefB67noFB+i7dGtAuQvx08RUc3+rpXYyL+o53KIugCtv
UBjeSx241NvlXDv+8VemKVB1z1J3yLnd1ps6tjgwjw2w4FJkJ85kq5GPy4a7jNzz
ayo/mmVw1d8syru3DQT1gKF7dGhml5yZepZblnmtuif9y2QL/rouhsdLb7DhT3PN
8XoRKtJs+812ElQKR6l1fLqy1Wv33+f9To0Pl2qNtPGiWhXAGJGIEG0gaYg7nyya
s+U9GDxyhceRhIXfjtNkBRVtDUBTxet5hArs9KpE2m8/JIa36xoMqs4l8Z3PQep9
Xhen1Ka55/ea4X3o7o0qQ7OSiWExnq2tGaDmzPzB7qh4Zmw0DkBZLSRwLypBFJnA
IOhpXViZWgWFci9X52XVNrmLS8N3xeOO6Rh22SvFiPhOB99GLeZ9ionnIuzQQMyz
3W1YrGnNAFXKacDULqW1MxexvS2et/DkQ3UKbyIDrdyIfxzeQrCbG1gopz0KTaud
YCDnaR0gPU9WVAQ9Xn0sfu9ultFAE2MWz3D6Mdeek+a1VD2jU2b7axYgePcG0y7+
uW7oCCStOhDXG2boH+l113kg1oy4+yIF1iYqyccb0fYfAx/3z+hDO98ecINwOq4j
x+LrCzkb70ZgST+ggjWM/6DH6j82YoyLKGK2XvmwKKzJCJ0GSzl0D9XYsCm0dvM1
Mk28NJWACYD5I27sfeGA1GDJ/0QAuoay030OIGwrafWGqU95jZZhQgVtA86uxibr
dejfaZIKhH2cEsedyfj65gpDx5ORKt4bXsRAawc/rV086ZWNyaJtnqnQBM6IVp+C
/PugqDXKJZHpSspbsUOdDJjd8YdKt26MyhBo6Preb0Javxq/5RBmhWQf4OxWgQPj
CzsnLLijWE3tqyUPCtKuWYQnp07ylQ/fmHCxMc3R712yl1xeNbQ+VqPxgmMgE9p1
twYC6tT4NYs7dSfO0khuSZpfIksjU6Ia+lDblpyLtx0TOagDbXngmKCULWftXo5H
4zvc6v/5EyGnC5hupGNAG2OViBFpQBk+3W2KXO8ug+0UbOtNn9q9IDtZ1bjfWAiH
XVM2WPRBdqxeL7PutzqgzQfzu3AHH3EbVy6TH3bDv86ueKrqaBE1E27Zi92v8Pbr
LjS9DypkBHnUpR0kC4V3weoLIXc3lyjIwFOw6K2P3WZdpUFMa2nXgz+tno/lSl1q
Owt9mc9BzBLegqXkFaeVVdARZO68dgVQ1tjZHwB78t+zV5Uso/st7r09W2T9dkqi
vrelWEJhHlwmgNMzAJkoCWkR6Mbv4D9wQra9WOBS0xiEQzAEHakRVC5d1e1cuZ2I
qly8q/T4FbrHrKcvk7ZEhNoEk4itid+ZnBeiu01YDx/aaWp9nK++ONWWfMrtbO4i
y5MHOYfBXu6VN6zeE3pcn/5+ifZbwFqW5IOvdzR0aa757m/nLNSxQ5O0qUSKLlPC
rbxHcqSuiO7hRwtN7nWFf4PlYRqoTT3kKAvkfKAejSolftIT+o6b5arnpC/rV/5e
eq8egbxCj4FDOYSruvkEd9Zc9IkScX2+4WJ6GitHVLDKl4fIcMqtmkOHeX6PD+fs
ZKa2HEahDesEK3BlZZxbnHJtT0QsI5wb+Ue2CyY4bc2smlU4MQcaKVOHU2LUAglR
gVXjyIWMHFFyUeme7rTTnaVG+ANJ//wZGeg47wtdFkWYr8dWhU+4Y8WdQ16qK1ge
QN+78kHsRKxMLMpoFRWK+KyTHhtOl0BTVqR8hpDhszA4xNyO3IWDOkPAMLhO4nJ/
NRpx4DCaafYYYNnTmuEXUYegcMUX4MTZ4/QDDDFTCzJf7i7YJhcLqNcyrBWgVdV+
ToDJbgVOa+8LAbP4phOxmnAvJpVRSVifEGVDqEVvlQoS4qAKO9W/1DPBrTENc5iN
F8xYuL02S2fJfYYtsLE2hiJhj2ZK4ZzsI50agwsieAU0v7C2v9uWvYOyWi/Fj8RK
v9+bJxMHJ55UBpCezei4Viu8R07K4gVpKhaAeOx+N8rHzUcZTltC/AjpX+jwEb63
3xADSnvulxFMLznWR5DQ/S14NtmfSt7uy3EdX3hpgMM51qeYDZkupnil+e7noqu7
Csusjjuww9BSqT2+YXeV5ghhuLmDd1d+gSnLbZ1dXh5gxOTOgcgPMcd1xH2dQzkV
PR4XkEM9FmhlV+Nje+EldaAlRNWg/VTVlX/+21nuFvdeHOsGdVnAewD4O/YG0ZEM
z+h+HwK95MRN/5dTFAbH44JaHN4v+e7jonKXiuoe0cB8xYJ9Ndeej+4+yqeCdA5D
QIaA/rUzMuaDT1knBykTHRtmgor18YLELo//HQCBZ1J0YxRfzYZZOXRqu4DytxJe
4Gsc6awDDUg+9caa0VRdMVOZ5+PlVTeGkt8BAS1RhwThk7w+naJ/Y1R/RoUiYUJO
dqZFv8MB1/h98MEBOVJ8uKhBEE0yDw81zVBsYQm3e+Gc9fLvBAGSApp1TnvloE0S
ZNYN0jFJV1FtDjKRZUlopN4Z+qkANPQ7Ig6pPfFevX5GRcrbt/p8ZDabsTweXuVx
sRuuszDgJHaRNFAIq0FFtmFLQ2cpu2w0WTv0AJ5EOQICAYQvyZ8RI7HFP27qn5xM
DJ2884r8j9ReIBq1HBFNh9YzV7Kc4Wb8vaEkLy/UW1f6ZPe6qBgju6MeBF+TTZD2
VgGt0TuWbnPlVbb3GJCjrXD77KslywxghEg3IM3XmNWTWmKmrY9wHVI1G/LMV347
IIpkPE/pN76MzZDf9mCQyMlvOFAjlHgzdf/GCMM8BhQ3CO7R4K/Eeg+EjB8V9+EI
uK8HfoFlB8+vBEg886SU9QjWvSfmwORLDZcz8x+cPIEdIa4F5aM6+7q/yI+62/zG
iCaMuPbJPbAhPsPtlK9vfWfGo1kSoPIGd9ZewMNSlkymZEICTfQ1rJe1AQiZqHpL
P5I8s22bwgw1Hn8sySR2gFu2Ateu3fVFumQeBU45bL0fATkfQLZuKQS1mgSZpy6L
aBDhYgAnyrAvE17vGkugAM1CwGFCgasJtMwv4zMB59G7yYOIZ98ipDkELb7idqnt
7Wra3IeQGSrwpGRI7TU/wlC4uCYyfww9/wYmv7h4k1ld+ZA9ux4Wyq0Lz7EBuabE
Cstmf3BTCEUVNlPdbp2t0BSzeba8zgKNAWb7QAXS0PYS6ldpgMwSsBi+qRWJ3XBU
NiVDzr176jmJGLWzqs7U5Qgx4MpSSNT7xIj5Umw/rwJ3pDZxInjSWXNNhjub8Ldz
MVUe2jxbpF5dtKYE1rusoD+0LWxHIvrSsud92QRxg1tZcmk7EQ+MWYQdjuVpMv1g
4fjqXnlt+83C/vIOh6VgYGwH5I9GKbC17R8T5aeWPCc0n95jWw+tZ0/16j1wnsyR
7Hg6idPC/GtESgkoo6Bt9UfIiBgNWTDpJIU/QCWmVtQ0kVjXgaNkMnIS28jHOLMf
Yo/1r6Cfooo3HVudgdeJEuhfe1y0pkPMXjPCpZJ70kXNEhu89VEpDUrPfm6Ac0oM
yoxpW3NoqVcK26C+SCSB1RW3+lCaYLzi05EknQwLQd+dcKs2hGuknThSaUF5WLMe
zoeZ+BrLmGS9fyT3PYScFDwNNc/4NIjdhvNWeG9a/KDMIYpDGlro6dKlQE7lccHO
0CyNI6iQcz2+WqDP3ByNfRVy6wgUu9lYZ4orkpQaAkG31IxTZYxNgRtt8+eXbLUZ
QUXyayPaLLfTSP6p80ACf6K4Nf8PqCWcNNdpqAWq6N5nfSSVhl6e6dKwwEJO2vs5
itah8m3ulf5lmkY67m9fTcuxWUyP2AOG6zp02mgqcbfFDAvxTuj3gXeTo7wrNcYH
Hwvdp0ERuXqY+AHNB0PYMJQWe60CC1PFH0S25TsWpUDcFCmvOQKDsnbOg+bgRkmc
Hjf0PAykkYsm0dVc44ruxgkQcygZKBsLKvbvctjHoTHAgZ+perT9rnvMixXRTn1o
CtiveVSv+LqTJ70VoYTi7zw+QOceFzwqvzZTSrgp66EskylQq3AfVBVJPeS6mavl
`protect end_protected
