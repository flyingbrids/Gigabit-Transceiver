`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
HbbFdeCk1IjfEanbNTngGQtT5HEo3ckC4Wvt2yk5sBHt2Ao1rvXc+a5MViuOlm9F
zH07WIUhl/QJ9f7+Scn0cGC/6NfpxNwrpoLQqiQv6pqLL3kyDJZNHuxbACa4Yfu5
FHlSvjIJYFEKS8Irw3cT14mSHCjklJnrTqMWwQae/w8ky/78eWG3se/4swGCakfn
ro98KkhY1k+oGow87soge47mQokTdv349tQTDqVFtWVjSw/xU4hgIAe4p1uOAfyZ
MRj9JqLG+vXbllY47vCy3JaabIbgo4mT43vxOJmKHpvwCrpH3hn7FB+kpQnCGrNa
xYU3Zd4lQvhY6/VqBY9yCA==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
LkrInqXO9QkfwjVk5TUb82uiY89J0JcOMJ6CLJWx/5Oege6KxrrJITBNxzxYYbuD
L97T/UNgq2Bt9C56q+bhw/dDNPA+Ng6uGGrjDE/bTbS94Vg+PCCBQ310GR55jalU
iP+yVZfQsd2xxDeKWFT3Y2n4Typ7VG65zdzKjUMnvFA=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 34272 )
`protect data_block
pOjXkqPVA1eP6G7l9GmbqQTX99psE5u/sSjPaOxddV/GyNeSHdk+QW/epUNmLNC0
Gpyk70/GyfNfzBzZZJJb/srhhpSLqIEvPWy4X0hvKDk7XLLQUqgXTE/sx24gNlDj
zbhtlI1RmsO98nND5EXl8tz+2Gnf+FazwlOyz8j5JVhoZepVBvgagSZJNO3OhP92
U+fx94pvz+DrznqcsFtgj03nAgPr/9ZjW7DC339JOsL4yWdC/O2G6eiUIZqIVgWx
j6qGBEaU/ajZCwZC97mqvpKFQd3wOvykCvonT1dBiWne3L6O9C9W5PetOyAXIANr
SUzhpDG5fh2ZPj5SNN/L10G9N/JrYkpCY+nniJgrpxd2+16YiK1eVFFT3hDxiJUj
nfDVrS3Sm2oUoNd5OlJhwhPL2f89MSrXWZEXnz/mG5YqUOYzZjmHXOu5oTF9S1vw
Pab/Y0dajmsjAiO6MVm1DU2XG8o9y5370l7yKm2swVQpq9zYTyY1jiwJXCxUA6Vz
MD9WXVDfT9VerYTSd467gVdp3jIge2IkxMGIgnlcBsH9RBwV6u/R7O0AsAGBc3yN
8KM4v9AhtLQkBTFlKUiRQ72dcKTTQAOviSbMvOyikPNLm6WmBNqlE5a4vJjwaQ+v
0t7kFwscuQ2Jh+CqedHikyzUGsu1uKXk6lQMA98DhE8RYswXby7Sw8hUrvwsOFul
rRcI7zaviMhMF4d8JvYnzk3oMPBDn/Jf1mFxwcC13XF3ZXWX2KtscQyokaivE0EF
DjGdVrs6MZWc8tWONv9mVzSjOArP6Fx+HlQNJ/v0K8PfIK2fwAQPkHnEFLp/MRUq
FFmTjpcC94rODtOtayYDsAGrYNcvMe2HcC1U14h5qI0K1ajWYg6I1CI2f4j6sIRj
E1Nfx3TmaiM2RyZDcGiNhlv2w14b0IVGlO+OG+pGzXLqHlVbD/JSfcN8i46ll2v3
6yicEj+sNHFUZYMpsXT6Jr0jeTRgmq+3AUawg2HZn3IvJbR3odp1bA5c+nO71kMC
iBiDWZ22fSnBZQwcPhJWMbI3U6mPfgY5jMA/KDCEHaVwGI6tsfkHwwX/5SErjZdI
sQeU4CdeJOm5h6owAPAKeqSYmwol7Cl+ztcMVVTd48H7gCM6Aq9jqpwifdx/nffe
GJb1vu+47aJhN2CJKFOcZsQciZSsPYb6PnXphzxatGGqpuk3ttUTKdeJmI2Tzs2/
kkvz+z0mY7nRRHrf2pu/qQF6eZQdtxxIuJMzNiAathLiiEGlZUHpfx7cz7RQh58H
59QmzmvOYU4DBQ38jMABa6Y9Rw4ntRsbSblil/2mt7sPHrRVVeLBv+2uKhn0uoOv
4B9AnLyYIz0dyeXVJ2ztlTItYc3cAchsDhM4x3kd1D+BJKFqytPtboE+Hy/pDtFA
c69l40gyRhFodJPxlV4NHoP71wi96jUtjPY18yGOnc/MMRLH2xdncwzGOQy8a8Ms
zh9A5Htu80/buqfbjVgTC8+8HswI07KgstG5VqCaZUV+H+ItHkKbCbvgFIS3tlgO
o3og/3H/R+JMnzZe1AktWf0PxD9DuoxpvCJWfZ3sNrwVHtxFZ22aperuLgf0mwWl
VrwxYJzo0X4Xgqtq8erNtIcpqPxYNgVrsaPFIjxldCUWWzHQjX0NhF/wMqPDGSM7
vh4uoeByCYXlZcdd5VJHrhRAFXmJhoYVRxCMp9eR0x2y44VURtNvxKXKkxWWL2vj
n9FonMkYHX0vDVu+MbbZYjavaQ29OPfCOn9+56mIgNKAuAfA0bRUP/lpnUUixXDm
/dnYKF67l88XllYLZCLD53IoCWieZ/nkFzaWb7ezS3xJD9YSicMdrgn8exLG75Vq
2wib6TAkpR15sWxmbuSRlti1NOdi+u9ogfjUFl6BhPNICkSviKtR4w+yi2LnXp/p
zDTTI6P1eCpHmOgppdo4oWlTUfoqUNtBXyYB7v3mFCC/ATPivxStyczxSWas227d
BzEP3rpRBcdo6rp+/wJ5aqeJKQl3Mb73V2Yid/nRnLYcmj01M1HwM75B7iI5Fmrs
g9UdlvE1Mg8aGNTnIQUQCmDNvIBzO4YiCvAe7UiUPaYwBsjRdnGv4DtpBNAQgeub
9X/9hSyHAoWTB2g3a14Ct5u6A6OlJOZ+1fpHdsFkjQOdHi3hiNQUkh9WuzgzHNLf
Z4GCxnapDjh+UjFjg4R07h7sffmk6VN4N4HEN2p6gs9hjdOzaVfvLsgq3e6X22NO
a4DqEd6Qclj1dlxqH1RFkrmXed9NcUUm1lPcQuk6qGyTMnWncW8MPUayjQS9J3nt
1e6lr9FW+JM1T7JWTZuFL8IkQ3btDaqIGEigk1RJmPUswyiEe2ieWLxaNuLjP+nv
YrDV0Z6sMeHaZCcvTrAB2joTbbxsIqGJNZPcrvmcMaBShHgvtOys/FwHR/tTKUac
mmTg3TICz543GR23CuRO38JVBXBcRUG6oUga5lBl/L+UpmmOludvDPbGb7srlMaH
g4Tq48g0cDth9vKb+8Tarp5WyEWwJF2qjAJyOC4g0rTJ2m/cvWHhKtjM2bf4kmLO
I9Fb/FpRArMri6HpM3F7i3lo+o2zaRA3wuHzcmyYhIudmto6XQviti4CBDYWBcsP
Rrx4U1qZMOLW2xW6E0TYvm9Zsc7cJa+3EqacwhKwrC+suwD8WsqDjBi7YbJuG/51
lG09LxFSKv46LYDwEQ1S3xYCTuAKhxN1V470JNZvmSerkTAQHFXYSgq5oZ0oAhrG
6TETXzQGoRES/LqNPmnh/NEZ9azzNOVEHv7t5qEn+kaY9IwPOSSRkV4Pzu1a3XqM
ygZi/rEh6ipNhlmvj9wm09QuFPc4Qbhc1ely9B0rdG+jCG1CIbyEzSZG1pQq4FIx
+qmUHV7/fxEhPs0qPeqYZfyEPTQWZ5tsXaBuQpsJccDBNsOOP+aTij0DZNmyh4WK
8TEfhLw3FlTdlW0BuMM8K32QkADpApycU8neRw2RmXe4MxpB5uT35GXHpm1xUw7F
vXOtijnl0L24P413OEgBobXilH5Z4pDMblHB0BkZswkRUczhJXWl/C5A8m8esY0f
jnsVUHhFM8HKlqqMbzPnGZqU0IvKPtzM+ZSzmUuqkshUDybh3gLp/pT2CsYthu0i
Q/vwpSzkuDwycKbruU8cXWpr7cY02sL65CdLbLSbPD6P+cpdoCrxUX+40po2thQA
EPQHGhIf/BKRAezmfIRjMK6PORG7QTY2BZtZpszaRLu0k9h6lBQ9AxXE/Xug5uuO
XRDkIe5v/8KjPyt3zVeeO28i2NdskK8h2NsUIwp0CU9MMntv2hI4fT0tCjSFdcT6
nHok25vfAiURKMlw5yuiSWIKCw3GrYkm/PXlkdD4YtwXPu3rbPabnEM1owjsnq3H
kIaoTAgXn7hg2bZDqkLZQCCJ088LMorr20xGqBRiCgF1G4E2t91Q1fe3ft7ZSS9H
wEJdykmF7F9GxAyC+zCc4avbXInW2lUjrAop8cojSd9oBpaD5pLfl6WjK1hNoaR9
iqAsAmLMkaIcBE0Re1teegRBAB0HERcN55soLC1cUY6XSGDAHgmY419pS45RIlZk
cA9hge2Q/5B3r56RiwMFT6AaK+16EgY+QkvrQ0DvLLtMRrhV0+fk9DiTPCXzEVKJ
Zfhgl4kIg4zBXmW9ZR2SHAlKjzqeA+RIpt2QWCa09P8VTYVhtc5A12wmYcpFgLq9
Uq3EJl+9uFvMEwpRKJXC9NDYxAsUuqX/M2UGM10XE4j1obTWxEg5lrrpjJ2NBTGK
u10jCGkpX7VER27N0bYic5G8i46B4A3yL4KGZAX0EYRSth0dxL/+5Pim8VVX4+Te
whw3GXW35SUc3wwpDkLGbqRtkXMYI4/QDKk12XA60jaW2vnKqtr92R82tsrW4kUJ
5NtXSedu4X4ZiN7URXKmXPwsl/JeGD8MT17/LOjYCG5NEHTReLA/ATiQKWF3Yiuz
fpc4SeZd6+kgpLfYhh93aTLFuhtSCw97jE8NHpDIuEXbcenCy5tmm53FErZlWD32
aUc5D/KmqKuf5nAPJArX8KOm5v0cFiF0FL9Zk50WxhzGrbDSDVkGmm4EqOj45TJD
M8crxZ5KwmdWLw/zizU/1AhGfp4ADLWzp+iDkZs+zdLljV1ZDJanCAjy7FEgFv2g
Zn5h1bQ9mULJ9zAMRSNlN3dfQSUihz7s13khIEQX4y4dP4hxOdlZO8yvS1nnjlWL
KY0hlZZ6YG6KuLGYheejVOxoWVckSiDolXukpgRyyZG1T8VjD20kYO4IvM7/+6Ot
OQjIcFtzs/hPtktL2kJs8CIyGli03FDOO4x1pTyaWuDieE/qPcUEVmA6/2ibgAeB
O1q3Oke90Ml4TrYEDOYnG+a3i0LZAfT0GHZKx+JVDwRWdxSDSexKRoAUhsTbLMeF
veLEjiqIseRIwwAVvYHx9LQF34BhZ0Rz7bk8fIRwzRUPWa3NydK6vABxPZnTY9dH
mRnpNsWNeOOGHHXgC9fHl5bB5FIMBwHwGErklycRaCfaW/BZN3gyH53pczWD0KP6
y4Frj3eqaryolEjkO2jEj2rsF2ehgMNuiVPpz5+VsE5JtwgErK1Rapq7Y1dlmzr+
89moS7JX5ZFvNwakHlVH5ywPVvnNUA5NmcnleLVuTTw4i/UopoLdJl2zWsOiMBFP
ejA7cfzjmCaksUmhKMh3BZ+KDtqRjUPliU1a2rfKDsILEVdA6KlXNE7vFgmXqnb1
KNCyKf7/51pZmEaP870mm4ZFSDongwrQEXwWvuIhqwtsX1QN8toN/MNHfT/ODDo9
YpPYHi5NPox+yesVNFtGjeoDrd7tEhvAqNvcVKJBPzItArmurX/H4pcQKWDrhHh2
pxj0M4vp8KiD1sdx95+rQV6mLvLn0+9EjXn0y4xi2ykAoNFVLvGkkQv7zJeEhheW
cmrkJeZ2Q8Rr8cDzLbs8ymKo/z6W4qwZTreFSrvYxIMkjpTDw+EsFUdIMwj4JdQf
7l/irzHsiKYo29MW63Y8AKlKr8jyAOW6JdS0tpepHCnuqLsMQgZQ+RMsxUzsNf6u
A+kVREg9yznosZwkWRUCXATS1J90FPgIqI9Nftl7DYAUUOSZLCVJZazldve1wz6s
OW39ZJRWDUK/ZGRaeAe9NCd5HipGzzKoTRJiBcxD2JvETTfcyDlK3Dirj0bTaDd4
tuJjETJmdmFilzG3ZH7jHeymCJbSC5Fca40jYPcG2EuGp0JKqqyHP/QQ3gXe6J7L
8UnSCqxkyeMb+3eKrvMiSBmd1q5zQX8Na3f8tnurnxfINLXIOfRTkKNia1XAQYs7
FIituZ8e171zIU+4mDSgncUHYgafRKBfW0AT7gCf5y7DLTgWxbtjdSCnr09BbJzM
rziIQ4IJuRdxage8xoOItrwRPOYhIROQX6o2IiGcAw6TIuV+BUXU8OHl8ygXGqIO
yCopsqd3zmfBuINSC503LKBQeKRNUMxi9OO+zelSaHfYZP7nnoLWT77ZdOYW3/n3
jFdXq9RUfO/cpgSSaUdWkFnd/fAoC6MRMFfd0ne9cPqywBMCQSO7DdCXUrpELNPQ
1poIssjLVZzUCdu/s9S0MdErAVxaknkpCRNNBJV7qBw/hTwS7SnVy3atZ8l+JEA1
074cDDX8NO/3Qt+/YN7rS53RxEbl2HhaAiZ1MMLNzXjpGtwjpHqKruAU+M4m4CVD
0thotHQLxa7tGzPAo4ZYoMZISDmbW7lEe2evNEOzZDp50FFcT8DJCjExqpz6M4av
AAUsOEhkL4L0wphwvh2xd6XzZYD33R79uxOPuAjHRkRkyO12d5zo9rmBwf1xg1mS
aHbeeVPe6BRSniNW7LheSEZF+mJ4qdNEOK5pFPicIMTTgI3BUZU5bdD8tP+yadna
XrOgzJJ0pRk0uoP8r5tRjLEGOQpnsy732aG3Ey5FaK84lHBD0wNlCp2SW3QB0r3Y
EKV9adH0ZWe0Hs1E2XLFYFkD+3hSxAp/2sUQvAlUohSv59htd4al3TfawctS2zQh
lrmQGr+Rg4/5Texhxd0Wz/BKddo3UOQ1GyuETRYsZE3Tb6vup7IoKeYgLMRZobHZ
QkzcqgKj2mktg+evtUpjwYDizxkha1MazEGdrQ3bVvDmsGPi4KDl3KieodiYrNnn
Jz3gPm1Ge+y5omGZpH3fSF44/OBn+tN9h2pRv4Df73KEnMYZEQn9uVAUEFFuGFgD
FP0SDaPY9am3xubLPohlNJbnsz/J/1+KngtZuOp3AEfNFw30WQms8BbvWCF+LleD
Zh0GRzSbTUfr1ecTOGwyMAUPrKI3B4ng3RIaWhk6OQusCGiCdBqm+wyWb2rJAmX3
QfKTfhsRCqzRvNsmQkDh74qmxbI+v1Oi0oIvgNO6y8logJ3gjYoNkRPOkzWpznbc
vGJHVWNdMPvhmQ8n31HfZjo8sML+Gy5dYKiYDrWWqGa2aOxDRjq1w9GG4Ow1R18y
FcYcZufAbXgUoX7tTzwH6BxguJAWvEITWdH5Rbo3EdegGCIOJM3EdIZbkBGD4U2l
M1ZAvYWZAf68Ef8XDRZ2ue8jGPQQr9HyZw0EV9h2zyUXUvotE0AGjfTtMF3/O+AY
x9qN/P+DyRpJbJnJj09b6chDj7RLAfYr94/LChLpTepwt3LAl7t/giomzq8NEQIX
D7+01SoDwWQIUtKpmtP65Qyf0ojR3wo6NJgrxEHHYMcCde/sPTr69+8mSX/r3Be6
3TEX6XpZ2yEpDAvEXcB+tH59VJ6FBerDQ0y0NGQ3ylnjLENqmiXTu//tOa0UssI3
XriQwpawvSAr4i0O2jyEnw+mSKCkk5JD4N9rm9ZLYl+cK4kA1sWnzTgP+AGoiP55
zuGW7W7IH84j+hYjMmXHWoXVAdhGignV1jYmgIPA179eIlGRbjMYY4KTZytVRPx5
qf7i5fymbY8e+qOrPpvSSD2R4y09FQyZ+rSWKRRpLjhO18Cgyb7yJhsyP9gu8Sji
XexTaYsc9r4rmNOqarJQbQMJav1s2pBNu5dauWkLYK9eEww/Zmfjc9E+5MHbpiWe
F85GA07/CTjj8qHTl2ZQUtX2ZpbfFpM9iHnC+DYUFtFSlCGw/nK7i7c11+ZMmrKT
E4sETpB/jZmUk+409QB4SaOVoWV2oRke8sHKD4wSsAjrn0td8thX8p1+b2Sd88On
YsYGubyyTKAia0KMuR1QqJDh9f4XCDSPU9bg3WCdPc1sC6jUGST9fyvcAiaqt2qb
RTvdRwDKN2EBnECc6QluR28HdFiMmWGpIm3VSqdD6MXc++cU+a2Iz4dXl3NCKtmb
U+xuKSWSHu+2CHF++f6CPq/d+YYDnrbfRbNoG2WXFTUSWzyb9Y4IUsm1wb3n34Ax
OWFMIDu5DjiuZaPk/iqM1hie3iUwM8ydeID2oBT9pVotJVAqTKqVtFRKOGft8fDL
Hqky5cLFkXqVA/I184/PFibUOfvvxIbO/CQzGKl2+wQkb5vGhrd858JTG+KD2HJP
dGVgnoFrel4Qk+l880IvFUgn7MSqJTWMCPmgrsk0Wah+hvbzEWqh0b89kW0FM21K
0d9y6AEh70FDNU2KA185g95tMPDrI6IAAJiQIPh+nIjxKT+Hkp/+qxXd+NoRYhKY
BFBHN/1ReVsqWmQutIVXCS/W9ZI/I15LXVMuJ9xzaWGDC9LnB73zJeab4X+aASr8
AMbaxahbzlZl8H6v0Fv77SiJpHguqeAyNhbR9umWy4g8EUayBUYNZ+5SVaI82zmI
GfyzO2+bVIPDrjpWc+F74Mw6DhuvYCOlpeKEgTjZ5x11MOD/bmdEe5qZM1gf0Xmy
Sv1h/TYXQ77hDJq1/zSqyBugQDIFlvPJCfqEVw/uhl/VmR8qpSnMTQyj3d9sy9Z+
j0ApJi2r5VJd1g4Vu2ck203RQs98LEFZc43+njedoHAepF4eeszfroGpMf6dDJF6
aDOU/fljUXOqUbMDT2WfoFTdx5OsAERabTGUt8KfC6mwYNqCvZRd1klsdjraqmZt
iniHkPFxF80XxbI+zsscJTb7zygXDCBeqOdOY17NREVdVVz3Rges85ufCixMb3Gv
brOAdVnyzewrVbySxSlX7XX89H/2G16Xah6r1tLgrDfw0EYYV2zampNzidCb4uGz
hfVhQLkBvQX8WpMVMXcqZaeE31vJsbhHBovRfpMQh7fzRm+J9MzgzcMXgQKY8UzB
uoynvxrrSU/mn5r3JcBL+GwbraFOzUc9uEWGOJTdNtM+2hOHIsYvMh4IX3BiWCyd
h63SOkFdvpvw/wErVkhL7aLGMcQ0H2sOA+nTpL2GnWQgLHQrW7kwVF0sEdfLThOz
MdUhM7UWdRDjy6L5yzthxfmlkVaVhJar8F4Wc9I3SEeFUmfmi5LYmmjlPCf54xrI
bqRzYw6LXF98n/syXZvuTC0IHg3S28CcAhVrKSZKPyzc50GaXPP+wH9fHvDGcG02
sVSEPjFPELqlQgSZhgWYWuL80o96wIum7XEZckISnooRZkqJip3NJqrbGJD1BBem
KHZVP9j5dKSzvS7BKRmtVCLWAYCeZ/UPXbe7JvAcT3DzWXFgxFebOm8KnEeess2L
jL4M/q6qJoFXj5GgX60wxf9/N+rT9mV1bMolgBKpnQip8/wkI5u6x8PAfsG0NNMV
m9xwKFU6JyYyML2zEcIpOxiyT/G0N2sCvO51Sdj9bbLw/tdjnlc0lLiGvZdfjJ31
vIJ74nmjbytuRTPKJq9B6+pu5AlFiwncicGuGaYVIH4EveTpjtIU/1+53eyJXp4G
Xrx3txAfmraFo8eDeAYMPIid/z59+T+IkaKU2zesLOozGZIWOoiq3a4xtRDdOSkU
IivTr5/OWZOJBahAYe8QjPXQqGYPqWZZvUo6WL0DO51Tza24XekiCzLHZGeZl3CP
6yC/BJmfN2sGuD6s4zbROQy2bK80w3LVehPraPPE0MJF1OmaKK/De0PUtu2zBKfB
IkOYq5MAyXrCmRLyYLkKRvORFSP3aHWlVJGsbFVCTCGQlgMNwUnR0oBLXe9cO20N
RDqy3LGFpODi3qKHb2+lTZkdVhGuZp00ZYB6us2Xahap6XTjsdeDocrUYvfhGkSM
1o1rvHbA4AWvvUiZDUWHzqd9PGxLVfvQPl75y4KWUfBAXY/D3OpScxyjuBwxQqGA
8pKvqG3UskYGDZ8jY/2n2dBBJPdh5jUrppnRRuxd8si4GTV7pVMDCJ5tyE+hRqBw
FtR0BQZD8hXlfeG2KV3eCEHjIcSkU7sAD84rgC/8TdJBuwkYs9anhkXEiJjSiu8I
ilhkp7QeBLLPrcY7hWeri/y1junnLgQPZRfReEnYv8LnI5yuFkKszXU+1k7JLnwS
6u2kONi4JmWpmXMTfgLtYtFv/hDz8RY1ex8R6HdIqy8QINe4tOi/qk5Q/e5IQonJ
FcVGC6oewkHxNCi6EuGbwdSIb2NkISn8Q61Om4qq61dTfeMiN/0xKXQI5E66pBEG
H0xAVnu+OdV1RUtEJxaRQEP1ly0fmxf02NCgTJh1+BJyfc23dXpRJuHmC6JBLZOA
u2P99Hejc1nuXayPGWAz87PwYNRdPbex8k4YjLOfOFXWYts7ZCh6a2pXH/Xs4sO7
NALxSWacJSzhuM85Kz8n/4N2v+cG1dpoqRtopaQvdpl+qSBJAS2qMuoHIz8Ml1r7
YJAqSLQcE8v6GxMi1JuEDVoBtyFdGGBu4BHq2ex6kp4THm1u8dx0E7DsvnNsH7Eq
gFWENbKYlUDC/JUC8TBipwNOgQ1qlNtTq6uIionHo8yndmzCUY9F2jRiPkSP3F21
PN5P785sEn1ZkgM5YLp0JDhR3xMPU4gSIKcgNOqzJ9lXaWKyXJiffz5tvCWpQAJq
iuv7WtXIylQccPfJYUVOp81uFcHNovi7HyN3Br71xunmdnXyqAUJUwaommrUZDoH
XMAnNRq2Lh5RLtBq4p9IhNlTgmxvQmDecGKDaX931NuV7DzG9DNoFTO57kMrYSdO
hu05CFsCI1oOBLZd+QFBj5zCBuSiXTxoTcRu0SN0O8CVK1K2D6mrjLn55kLmk7d+
R4RAHjLT+Xu1jHrurKg/Wcnq5Yqc2KVnwSXp1Buv5GDo20xs6xzmEVgqL0lJZ1Na
TvSLl2ZT/uEdHHnJF7CX9ILq9TtJVReW5OYR98EvSUU6YocnUzJz+EBw6zV8T97A
Dartog+op9KoHb29vi9UyXZo4ipT3C21RBtd0EPKpiH6ojNaiMJ9R4oCGLz0+Fhd
O1I5HzYP9CyqyLS5LyP0u0SFdZKFL4gy4tmAE055a5x6CReUTvdSqiG7E5aoSDRH
tzMoLUZNVx3I5nIvkDjPtBX5CatVcqFB7MfQLEgThWic+2RI5mrSHGSvw5OmYmSK
CJZOGEFBUpiKQU7GyewDiwmWXlTozHJ6FeWks7jN4ZLo3S3vdPEZml4YJGa/O5Pe
in7O48lHMzwdh7j/hy3UrnIynEaorywKemUSv5/QP4rupHKgSNoFH7ororgNKnSQ
t0rd1IkzsPunn9MYf9+B1GlKLFboZHObZvNc7bUmTsIAwZVLvJTXqoPTsUD8HlcP
S4Ia1SJItuni97GIjIKbbANS0be5Vp9oAleqmn+kmQ/cAzIYNLAOsrH+JAOcMX+n
Q5SUCNRjCHas+8u35/y0FwKHh+KEAeupu9rkPaoObG3r+6cKjCaQDUudfqQ8NKWU
cBuucrerns2NY6w97AiBUkBDa8PlMYBHA8+0gUQjC5qWnODG96E80klrAZFnN7Mj
lZ0hB6y+DT1Ocvq9FqZ/AWDLhiWtzGRqOnRuSkLjhKLGwxv0iSTWOmuMDeXZzwM+
sfxVTZPwKutlkuLQ/+etyhjVcw37Df+gRLojdSmV6n8bqJPaBMNz13VWIzM48u7p
FJkfIt2fH1PHiY7YszsDWwU+bzIx+/9bU8o+7b1DUbM1Rhve8n0bkzkHPTPKnq64
geVFimxLkbhLLUqDEEa7589AvCka62J9CAJ2hmbvUlB2xPGaUOjwOkUx29dFTN58
2M3n/ItV9SZWHGACd7gbWJJrdQCSmC0LRlobCHR7CLl5H2PYnhX4eSy50AkHyzu8
q6+VdCQBuIh+fHrGD+kV1u7o0fW9hxdxEl/vUGmdxkkdmUzMJqZvFM+jYm+m/U71
JCFcJSa96hj1iThFAwCdxNPo9hLwSZsei4mWzzdVvbSTw+LLH1i9CeL4OGvU+htK
LaohjF3FaiClg+JfSbcPQoDblcPL3XMJV6X7iEK37bEGspGgJs6QkdnxnUsf/MNw
mzL+srzZo/0M9W/V1S8jfSbH8LHGrdOJO7Zzc/8QVix5MB1HJ10BQ2Zyof3PptAW
CzIJDo+EVLpdJMNUxEpEAmcm1FmfUc0UVULsWmiT4PBVBpBuqNDevN+gvxKaN8ar
Dd5TpK+XfMhKUYQ4+Ig4d06hltBnxB9L9povFS86+f6iDEeJRBxC0z4wJbOzF1H1
JjE/MLdGmUgQS8CQu8Isiwn5eoSiNzhqcre4tkwdpRSgQapFDFZJ4iexDmC71By/
Aya8kExHDH3ILJml6cNu1QNqd1DuRcYFuOEpCAaKcUbua2uX2IDcaA3Esz5J8Ok4
7QfpKV2PAYu9EVFpKhDjaC7JmDd5rmJuqWh+owk4ouJiuuqTLktCcfdXfAXqzSWa
a/fzUfkkPRUXqxaC9H4g4toaidzKg6hBprqrKnL9qLqSF9FCVwHz68uhRwolizRD
Nwvbf9aJqQ/7GRz5AF1QXDzrfoVyS6aV0JjqOyXPr6wIXVIlEyxaNJUZzqF1qCX1
XoYirftitC4LpTh9ypujzMuJdjC7Ez4AzQAnRn+QF5CdXKuIAOKgEc66n+ZMN3Sn
sOlBhFgtrKuTK7WLWO6QBzLOhfP4294v0WAGdIa4bG87bnOaqGES4XqR1MJnvrhk
RCQMEtu6VpKf6Hq0w+kLkZsJRVrObz0hm+m3kInysDPf55X56H1T2Wyy35NTAef8
4RAGahmocMeBRAPloTfPKjx1Cv3RbnGwRZJ+dic/N8VafE3j2VsKeU7ernsYVzCz
bA7Y8aiI0rNYnfrwLcqg0pyYZfO3xA3UoMWkjVCSoJYyDJiM4FejBBh3zQcKdws2
asYNd53VhW3zjyAJokEMuWsvjkPpRTIOvRHzMXXZR67xPoPCmkFqALQGaCArRUkH
W/wcr3xoyRi7n6nM59qcmSSK9nUta5RpPXA/9RVUXl339swAqnelqE73howy8qKE
mHHncvlLvnqfAYWhcbuv+vOmEeljj+dUl9/jSaBru4KRZ4ZMIisHc8dH8MXBwGXZ
rTJZdYsYmL/CtsrhBMyk+c+iLr9G2BCdEtZUkeqjDXfG5njDeaiPK6/GWTIvJXDB
fkOk+ixo2PvZRpaO58YL/k2is4O0sJnoMPoAk2dDKRmbkV56tyAUN+nSK+HpSDXr
4fT+/WhtxVB3zRL9swrx0+RqECrtRj4VaJ75lkPEythR4RQsJwRrxhoXvi8N5x2k
60nvIBt/TFCvAiXCAi3u7bzUs12rrQmsDVFTvGnhdtnQmUVCXqx+d+u6KvcSJqie
8ZeNO4hI+LlSXNNbAxgnfw8yjZCuyD4/QlwPJNXmxg1UB0gp9biagZLqTBd337lG
RZI7+ulvwShtG57PW/Ci1y8pHKDLEP2aKbL/4xvsq9bcdULQ4qfqVHLBmybYo+Sy
8iG1+m9cPpny9U2kYQyxRb/q14Kc5BQuxT8bpEdNW1Ihxxpx46JoCv4kRweomVsr
PxB32DC5augS+Gz6Zgua6lavSE39Ve11Ib+J1N3TGjitaexTOxqooUOOhsnI2rLn
OYMOQ/F60mWkOm+9rDb/w+7ZOGBydcSA/ICT8YQWecKwguoO0z/yEvZc5diEWGMl
9L178ahIxFsboUfvrH09bc/XNMUsv1sSBGHSxF71gSnWuKg5RaMWOC+WE1dHJwLK
bDORMSZSvc8KupNNTUH/QEe4dx4aMCFshQf27uywV3uL1VJ0Hmt4RO5d222bhBQB
XzVsNWqlecVSAWo4Ja+fkaJJjDPpTFRw2CggkV82a44ox+A4uruMqlBAfxhShBo8
HQyr9ogLwISejbVSyJnc3AyV5PlQQiwYVYiROwqGj9l1U5sR37alnZnx8+FhZVFk
9FHFbC7VPvt4ME6n9XdWRBCTUrRRFPlRDFdAABAikwPiqnfKPPD4tTVk4TZBJn9x
hJqIc6Fy5CFOEiOGlfFgmMCOkaChzg7rtF7OX5wrbtjB+oqU4NTIYnL2Z+SchXg9
aGT+TViDywRGG1oePYbW81iJjPhQXk6MhLxV8L6R4eVeXc0pkmQa3i12MQsPNXIW
9uGbhW32fnLlhQA7FongCZ1GiuyupUACAByFN0D3y6P1oySaYi8hshjh+z32jstk
6ofLNEJuWIsEMnKDVgZK3KF98rknTJV2xOUxXLOfVAjTVFbitqBWEMU2YnMaYXP8
Weti6gsZxRUA7NtxnzSr5ad9sKRqqsEBl3IFbLoomvx0v9NNPkqDxejZDp6KEOOm
a6b0Z3wX35872NEkMdH6mVrJrEeGJimjaRcjE8RQecQ7EF7+VO2uKoUC7tnD5iD4
uyPnPY6bOOjc+gX8lP2AEBuQHuqJnv1SFceP0qm/7aF4id3ZJfXjDfQbKv045L5B
U5UrhMs4s+3mZO3ZH5ZOM7Rb4OM+dgGGgQfB9Z+21cn+1JzA7Tgsxkq/R0Wlo2SH
C+bWTXk3PgUdTlCO9o+Q/wMkVhq/OObLHNgpEcbxUruhBWtusqlPbb+lcEmOyJdS
s3jKsQmggAUaCE3/jE1SeOxf6zHa/xN7Xrtu1bqjVBZKXvhV9QLCrfYEfpUstiLf
83mIRS59SUwFjaFBEXCC/Kzsk9BrcP3wdh1D9PzXVtJdO8WwGOEuNFCQdIKyFGU4
4xOrNFSdRunOznzwVtFexl+/PSLTY0EExtWkasSqmEONvcY+O6JPdHw7mhs7/PFI
NHo4+DeOdZfWyaT+8pc56IHLsnMheEGCADiBnspZ787YIrCra8Hj6qJ+gC69gcuO
vNIrURq/NBQhUnyCF4dnjS/a4aSpg+calrLbiEarIF80nFO2pVoVmg/BajjyfXLj
ISEDF2WD+wkz6EO2riLR+eCzKzPxpL6oYTCZauJ6/9DqCxtYpqCqq0LvOn+LVweB
PcQsGXS/VGiwpOPL17grUjAVb9dKuDu0ukV300QpDFXhPJPvfoYAuKh5dGs8Z8Jp
3lFyO1ZoE6jbpRwsWqwST3tN67sdAxIFUkMK2gtxKSTEVwmZT4CXuxwpysltyVYN
0rxtwy4AETnEbr5LRtHk4nQ/+82pPRXDgpPwlmyDw+JFN00d23/5wpPv1QezAStI
32rsgGCaCXlR9pGJ7qIOpb/kTQNQluh4qtRmzTjUtbCkzVqp0SzBNA241oRhDD4R
zSDL53hsmk3ytx8y0X0HyeQwf+En77L9XgUFSCUKymswwxWwoMgAw+hw5i+JlGAt
5RueNQ2tcHFag07OyK9TB+roxRpFvhpf+q8IZ/qYF17mfGgPAqR4Q0yFpREb0ACm
N1ma1IyVKQfY1IfqRf8MqFDvnbptoXeTFrU1dF5chOBiFFqeKXhthp048cU5p3UX
t8zxotsmUunqVw2AR8DGZOp4vjtvUicbPEde/FtxO2ASlSI9Vg8BQEykXHHqCudN
ozloHyOtaGdxWT5qFM0l0cM+DWd14YMdKkf7jgGFwaNUs7XpshxOW1jtQs4XxIk0
09/bNME/x10g5vvycKiU3Vzg0mVT9aoKWPLZTRTzyobA8LTxgq6/LJM813RsTjIi
S1HR42FJMAvRsklEE5CMmV+9ZRv2pMQ8v4NZeptlj5tqsjIfC2VLTJbiDmEF/DQA
vWHEosdxyqlyYuper0o2CI9aoSrVphPBe4eExbKkWN8PWd+qpAHwUHJCeu2l5lfW
iwL/U2hU+jhSJyqRW8MbFZRfgnbh5R6ES/1LQLakoZEhZapPmKmG7d8YAX8QJmVg
hH6aR/i7YHQurYQ8EbSQws6v1YEux1U7LCC6uzc1wKYoXVimN9akQHsXGA+XVUSp
gMyOaPAG1s253PjR1xdrNAJWDGqYfLz7ARozWVaqfefS2YBtyLxO1wUB/0qDLQmh
k5lRcOuKc6duHB50tnwwRFs7cQLYGhYllNeX0N/GfP7vKAkQ3+cv8I5XvT/RR8on
SGskbd+a00WXo0HGubZQx/hVQT04SthEwRukjYe4kwvbrJ3hQyfbrUUhLMdjSFi1
BuZv4Efkh8ajTnIxnDGkmEJu/GRILdsMUDkik953wJBlURMLkBWlnhjbcUmgpyy0
pmNsa+h3fZxKLPD/TA7MVqfCjgS1HwT7dn/HR0mX1m+MEvyobN2DZWBxHQRDc/Ke
l4qnojNiWPu6NDmpKa2gauT0ri+Tq6lGtxTpmcUGxel7r2JnmY9GWbPUzlSxHH8S
CUpNeDhAFvBkUUNCHbfXF+wP5R5zFDU6fO7hGfjFoKKpLm1isA2tM2KWV+VlqOba
JrVqPe2SGaktDeexVWjnCUvfZEyGvirDcTTtoTO2cJC3ZgF1Ac6aNpDLfOPZpeDH
Jls1zOG2QYJ8olNYMvUb7PbdF9meW9eiufCj1ZjiN1QNCPVIq1aRR8MX2W58F0U5
ykcJO1xsa5MsoAD/AEt2qf1eO8X2ThsFL16KrilyQyl45TjZuILx3iIr7eN7tkGP
vCS99TKnVTEwiD9px9fhUCiSjq6nJyvMOBqNFOgp9mXv80y3H+qP4+NOLLmZlipd
qrsc4BUoqYNE7OVm7jJWXHLGTnuconhYzlJiCnSMR9JAzMlT7wKJrQQi8+xlAhyr
frmoxfLKBrVyf6iSBR0haC2Uk9veXl5LCCypwTbtbtKGwER+/JD3WMNbxeurHaCo
18GxkX6kfDGJ2AHu/RFdOO2PlXFt1zHLTwaOUt0q8IF+SITzM6lw5dNVf0tOPDsz
G/n0Y2a2tQsumi8VFLmOGeFYU6go+1fc+YufE3rsFbM8pYOTCrvaV/Ahy/CPrcYq
59wI+xOBdxNrqL/UBHdDUc87L9WiwEFgslrEDqTlKQ+ArsvvRNTAY2xxLTq6QHJq
9EtSlxNdwnrC4iqk+u+Eq/6HlqM41UHwdtbsEWs/nL5VX9oVb1cMdp3lezcg10ED
LlzVgHok0AqWuSUp10cuqc2EeGvppyGtfIz9MqQmhU2Rvtd8sf7JFWbnRm0wnNih
dgqYY6IhOozPIdfDToCun/YDyL7CAzMopi0xSR84fMIqGmsL2KjoCoGjmkAPMZvb
vaobNKRNNGLNjRX0VDSfKSelyZkmbi5G84SlKzIbdYF4JLBLFfgTh2JyiCetycCg
T8G7R2Mnp8fDs8qVIjy//XcqJ1gRjGjNDawqEc+Yud05CqdFLYw8MEPnbbUgBBeO
nRapgpfzjjyyljYd/0cr0yhEUrjpE3S5t68ivROCuegnZ8cCldBiJvnfBZ3oncw7
8+YxYAG7QAMrgLaZ/JoEeJ6K+Ai7EYBO3vzUc2swcOHxyOMdckFrrnPmvHQgMPIL
KQJiHh1Q1ypcpxWKuH8W51uITdk2uE7Cf+GeM68q6FerjJbzQKyrIDtCMI6mPUzE
NJKye+D0u7SBEpUQBuRIxS4YSlRR+En/k0chnQ3e6MgBMfzmaTYTfrmHtpumaEqs
YW5yBNESc3Hos+6GDdY6z+4pLbLzaPUFQyF8C5cbB94CSSa3I2ePACGaBmn7T7D0
Jdhuy+moiMBGzba9KuoharMYizwt9jqPshWVxmkrV2DxtFOZDlqhUHyhsl1ys4EE
UmTb4wDRtm8UaBL0ijncdGta4d/OPj9CaaP5oL1vJ6xPQ6Sk7jmjD+dDe032xttM
xFSg60s42cUjD2PmnO/uGeVWkq0jcEecluj2tJDBLgY0WNglM2yqDcwQLWs8sZCo
KZ4TbmqGXJ2zZje0GE1RvFUMlGbVNSwbW09E3+wZLafgTyXN1yAhoMN8mvUY8enu
384kERJHJVzm/U1CSHH/Ptg/Ln43Q0MTrRHKKgc2/Fkrq6Ese8QF62yD7M2IbwrD
PGdGTvUBT33aT4zjCX8VWfWVAc9xchNG55kJCYo7TEYyNYtJK919ilOex5VIBHiz
wirlS8POza1omK64WGJJ9yfWEyhRrN9ryGWvUeMcSf/MjIUxRwRp6NM8kzG/5si7
bUjqJ++OO7gP7EIlEHqI9eijNeIBxtxGAL6miTkEIbYi60BdV38ka8rVigMVej1W
09++pJ0nxoiYbUiVBiB/LrfsvFIdbVpwZ9BrJZySfCm37DYkjyohlT57hFxRuiFr
j7/ySWMmxMN8Gc9iTbQtUCQT+JYKdie9FYI13/Fur2ADNIp4AK8tmmripQQ8J1xM
FRFdjoSBJ7+r+OS6EFegVaCzNWug5K+kX5YYeLbiyBMpLSlVsOCvxSoTznxQfxgK
ZksaGHavRGQFw6kFQBaiHEfbC88HxzvONO5fQI6wzNbRfHKDGVlOtyP1M09vnjFn
u9DZAfSH1sW4xj+r1z9W0mV8UUGW9T2sS3hxVbvY+PRlmfsQIqSidUcMeAaGv+Mk
tawstJ2xX77NsYXFMGd7ywwhxwBzokeht/aO/6Ewbq95U1WWHj0JCLJ1XqEiK4Kz
PK1vDAlhbzqt90oM3UMG94PM/uyu0op3X+WNI0qsfiaqWPQAGFlQi3iyGlwcLZVj
lE/1lUU1hhCqPX560NlLovuktkzV8ceVVyCCv0hewlajO3NUuwh5ZdX1B2YlgTl/
qgXQ7DMqycDwP/W0OvV26Jc3lrFPvKPmpiy0cdB+2UfNWmMu4Kl5hjNfCG3E/+bE
TLoT+HZeBLWDbKnSkPCS8E73eXNEsA+Hqw35htuZaYQBrftJo4/op29A3mfbb3Yg
NJBAi9eAZzNo77TSKtLaUK0dGSajjnAHoZXeTlMtawHuMUkB0fTz3Wb8539DNYEU
d0EsE7hd81rW2WyEg4B0bzyA56IV8Sb3JqAYxvZn/r3plY/FMibVleGnNXgr4Q8i
j+Lc/6vI+E+bwZTbh/DnmnOXctAx0u9K72cBYyi4RcCuDZKzGPOp+wBIMAkcL/7k
dOSaRoim06wsws4DJcJoK0NiYZf14mlq+GXOLcIS3bIjbOVEE5q0vCDucfwz5/3q
KqPm8Ai3oPl42if0/jP5bUvcsVF7sDQb3VlMFNiDzEUehuA+a29YVp9F/SYLpro8
3sgWAXsMf80KgvTjTFAyqrCKQzcvipPWvSTWg9FCqWhi2IFssBOvzs9EjEPgIApv
lB+Q3/vAJ64uHu7v3tH2DtOPP7cqrHmW19fiOzKZNckcorleVAb8QVs1Kr8Q896E
nSpHtxGHej/54ydCXb35ttZ0JSPUTxcnfSds343RJ+ZQDJzZS+tD9A2ThWuEgW05
IZLelTRdguiWNcJEHPrBYoX+nCtDFqLMjpJ8t85BvCJEnA5aqObgbqAvHpjIlL3j
G706ZE8UZ3ZBSkXzNq2M8M3sWjpLoBf0A0FD/GTzArDnBvURAqcRL80h7tAd9QgN
R6ZS3J61zmipY8WTIwBYeRSEf39z+B57UgQ2+n+UCr0m6l7SgIiC3ZpzGa4pEft0
WdVUTVOwDlxeI71+yMMcmuRxmYDLwHUMuj9cw9q6w/mAghpAe+OIjncTQ+JGf6pG
BvIjqQihiloGKo1X2msh+uxFSilXo6gdlWDB53+COdTRGQlUNgXRUZCNpG9tuxB8
sRaaykQIsgetJy3ZZs3CVpk5tDlEpE4khe8Rjl3UruCmalLm9DVhMSBqOkmMuAcU
QlIYHHNKgGdUOGJZqgUWtloyJ/6q7aCZXnJphFRqkaDE0p5RA2I1icY/P0Zvk8nS
zjPBtzD1M0q0fkiXjHmXJLYNbLMAvaCguw11NN9/P+ANhWOxs5sg785TJxKz+AJS
RHxW4TvdJwMp4tOcpFtWvwWod9EfXo7x+LIJcf6oGf1tke5c1bEDGIawYMTjnBNM
9q+RJ1U6oKPUo44RI6gC4fAyUewKR8TrPU+Uw+1+11LCH+7rtlcm3K8pMjk8yyYv
2W8aO2MPRPrGvR3ojV+Eh8uRbxNk92nyT49sux0g4xm7YORAls/Bns0DGetWDKWE
gTmaVwDsdks4E9ZZDbyjf/GasviSg2kU6v4SIYuteUeOYVfjmf/ZyXULh9MBhErY
enZjNbWAZc7djWcKBKfHvoPpssjrAwCMC+R9zXkVgVo5oDyJgXbKbLhotz4xZmiz
O2ry9Oc68lCBFHw01O9RMiAKj2DDjiWO6pBuXYvMIJENA0fnMsbdGxVLH3WhYFIm
Rr1/+YLgjsNmfRQ5kd1EgxGUx1Fqi24Jtel3fjdQcF9yUHGEkA2Fx/qHwNHaTiwa
mXJYsM2d4Jt2sPemvej3uM1Hdj+q1leYY23clAv3czG+Lsz2HjolNSj5edroAolu
AsU0ZM9z3Iq3Z15/JFZrBRpxnAFn+5xoOJjkSVUej7tLFq1kLVAcXoZWxsv7GBdK
uQIF02Eh61EaPEMK5dgjm00ibN/wB7w1C2NT3wRyACkq0lS7PCh+x+Yg7hqXfKJ9
fX0XdqJBv1t5mU+UioUSF3oHQv7QQkQJNO8JZtX+3rvEUnFaKvBG4mmPlrXzfYP4
/64aMjcBrsUjtdme0KExD5uS9jBbX5H2HWET6naednbmFjdnrih37R2IAU8MTHjK
Yqslt876I2WrCqXL4Jat2y7NEiBb+XasrXLgGpRTIt1i/QWb4Y2s9MrjKwx3gqTu
DS6Vv7ukFnkSKOUQO1KbXEroSzbdY3VOtrwGQ8ZtL9g6CAaj6c/fTEzbKDx2eh1q
SRJOcu1Z/ftuo/oMfSgna3fJ/rMc7VmhtJw16tCJFjDuUr2nrCVKNGQZCmGbjpoU
oV705WtwOOWnV9IAMVyvPDFgp6eG/G76BZ8MDIFOq/n1jzIeZEXDZzopaydCDokn
Qq5wn0rx/uXhU5VCbdZW1s9G1iVHLzm9XyvcUG3j55dEkssqyHuu9pyM67JgJyHG
M/mwj6+i2WzIItp+104YZnNA5+u0+f4sxiB5aSgR45eyoeUMN8pnE3OhBlW301Hg
lmH43vv3/E1jeFfAUUHPErbu67DqSb8rC42/+qSWtZ77q6BVMdKRVmxUnXTW/6jK
Mf5cL9RgLOP2t0jCf45gV+9Z0OTGQIlEsjGLf8mtQR2etxzgkpi+6VTT9H2kQpYp
twrjWBpNqV2qND2L8X8GvTYDSGmPAMgV5uiZA4TX4sc124nZ19XMqyJmmHdmK3yF
WdQEmO3bSTApr7xyfSNUkIgE8ltxXh6ug3HSX5KGeHJ5lC7trr39ZujB9Fq7k7I2
fpPKviYHWKlyptxLQIZcoNIp6cN4U92Palhz2N/PcXcSZc2/SsjlGy1D75VDseM8
DapGrK8TdAsNZQPoeJUXgOk37956Sme4sSGCzdCFPb1GTimKjQMPyWSQBvCAJACY
kxoi6ga/8vwEn6RYWmJcalbjvckGjkmlCSof68D50U8KyKrwCZIEd8wgoNRTE5b5
A2MYhrk1XoxgO4nBy2vYQayA1sHa/2/kmpdL/vmJ1QedklrSTHvYTyksIKGgY6U2
eeCcmd4HkuxhZgk8jGEXBQbEi3g774nkcojGJ1XHhS4WYUc5MdDwBz0obhbqZYrr
tJSSKeAYO5Eqxl3Wr2GW6j7boKDD0bh+Mj7dLoBUsvuwlaBuCkwFQTH3SoLzan7V
O/PpZufFSOORNNC/q9z7t47qknBa7tZJ8MaBYOeDZXn+LzI6N0Nag+CkeMJfCeSN
9f+Eo0HnOHeba9iaWNX5GALoIu36Z3ZQCj/SYmuSmRmnbz0tmToJgBVAW3SgM2fa
ExBm6iPbK31mJvVv6HSqbMcQnXIYKDGbbJ8Gy+2IVPhTfjZuoxQv9uuBmflAvs/v
7W4Yw59f8x6eLNy0XA1x02MvFJoN3HNT1xb/T2MFvo3gow+NWZ46PW/c066Inl/c
tEUswN8fgvJxgTdao68ihjVx11EH3xakEDSgS35IYosSYMmqkg/SZsS6lgM+H4aF
oMgF2JN/2rqxgLSvVfljb99Zu4WWnV3fpbXyV0E/3JWqoJqfpaUwkFioMZPk7SnI
oAnsZPLpMl9SqrohCbw4aqQSS0A7RTUdT7E+/Eq7llhdGxNDbKQDwKd5XS4ipvBQ
0mY5qm/tSPtjH98xuVqhm/n71R4XBSO+gAz9DS4CDknkB9YiFSq1V0+Ohfzf/F9P
5C4LEw677/Ebj1q3KTWfyGLuFIPpU5e+yRagnmPa8ZzVIfUizKcvCrqmsMJ9xGef
dQGdNRCxjZQaqF0ByFi0uPDePteDmnScchjre6wpQwcMujKNqjuBDv058wxv0ebC
50vfYVr+pgUC7mMr2eYssA0GrjTnNaFJb9SXGrO2f1Rt7wmqcKni0zf4QGe4J2bE
RHDI5d6Kj5IvWm7x6hH5tXI332hFyssK3BBTov+8+2DF1EKQEYJnkcVmNinmdSN4
vnv/A6NiAqgwI6Xpg5xsXvpL+vTt6R0VIITPgwc0E0fjPDnFWTEAj4sMgXQfVtw3
bz7pha0yc39DrWSaskQLmsYnm+DwuCnKfi0Yqve00chXd7bKOBGfUpmfZ04LLH6r
0/G6vfXM/CWWJeWTzGl3xfCAkz902j5tDLfbWxZ8bhI0d2Ok35KVoBGpslxPfnjx
apAB3SnRx40pLjapTElhGAVKgcQUdSJFiDxCABe8sapPKxYaLQUVXIavWDjq2Fwt
fRoc40EG+Gc20BnbQf6fJo3S+VIzlkotRae8nd/QSCXM6Vnpr2OSmBXgobhU1Kar
jGK3Z/J5C9dPu7nevTgqP1i6xdF7yJkJ5kXRPM9qIo1ZunMEkVrNn+k+Kg7gv8yG
DHzvmBwuxOk25RVihFYUUCbVCKpg5Bm9OpXttQh3ere1dQmO/5xO65chSUOOM2mC
aGH9ET2jz9cP8EOShIy/K6bijp5T6CLEyssqmPIcct2ojXm6i2FyGqqMCz2bVxiW
S2HHQYn8AvRaTNgUwn+nNlL8nmhl1xYvO59fKRxWfZaHxIpNvcdLw6kW03JQmtm5
uq+UWpnnL23CYy8yfOTsqAPnMO6tw006FM5hg6MLimfPgg8klw4pMOXO2yn4P3E7
utNA/uOTNbC5UuQuLz7RHKOHkt/3O44+MKr3qpM3Pv+vK3jUV9ewNkRKLa7JgD91
ricG22WQxFMvzonTpE2sCAHifU/CrKptp23WFdNSJrQnCyFwYIvU5PGvLYCnEgCg
wt3CM2+pOsHmS0GThUIOpY7p5HGXJn0h4K0mEzWbVffY1UQk0De3nsAagqspaWmg
JhYZLCXan2s5v7q9QX361KE9SQXX+/r0hCwPZWxVOJk3BqrEB3QU3s+8mNvaOOlK
vcXWdIeLGfd4RTkdwctKByQgcGnd510vgA7Vv1LvVky1QUrX5Sd6mJBZdxAWMSFL
ukbrfzNzPboWvayqbX1V1FQqINARThlP52i6PU5Cqwz0lGZ5YupOstPAApTsn1r6
XPmAtYqcpe1OCT7rRkqDFqn4QRzTDuolXGW+s6GH5Bj5mevi+9ggI383MhlXt7iQ
uL8nfFLS5q8/MaP9BkAyWA/BnjCGGHJ3znkcGXv3wMffM/dsXvmususPhp3mGD/W
9QlNkcyxuCWQtKcURBAWsFFR2pRGdz0j8m5CcluTwV3zBqKolUbKCZUsgJvW52PQ
F4QeneQ8neqP5ot7ZIjcsKph0KpPZuns0txjaGqoukb1t2Mjcdwl43w1V/taDuXM
RUaLM+IlK1tA9dh2LmuzSuM6p3M/pNLBj5rMwPJ9FMqAv+p9zlyZAmEpYp7HonA0
nyyldvdWb8rlO/WQSns6dlotT8PmoXzbpoZ7MgVessEJqXIac+5JBWsB7vL8V7wU
ixBhw0O24GzlOXUrRXC8tOnZ3P05mkciViK/Lex6CCdDiP7mUgY+tljryUJwQG5L
/1bMhzZ8BUkx7o6hLeBdzAvKRCpFn1jFxxNKjpqHqXuEykCPC6ov/WIcqL72qVo+
kWO6lhF3tacOyuCGyHGzmGQomVc05WxUyD04tb8iljALmjgSp6Ecv/r49Tyabq5n
X2FdppI4niRBUKLVf5BQPGe0WMIAHrBIkALmSwr8OZwC8MLsI7d4I7vW0ZfDYSzm
74GZYxELxLjSG2b1EcwOt+qy92rqSeFE62o3PYecmrrjJnG7ZznjXo+5MCeqGZfw
7nyoWS71oB9Jt0SFz07uIj8nQDQG5eiFzF53m7naB1e/9X5vND2E4C4cPWatSFQr
AsYexeky6ZsjvhCFhWIexartI/eGfFcV5SL3s3mvjc5Ri2FbunCHyGgHLrX5wJBr
k49g4S9h0MIehyFXivhcUhdIDbVL5TlLfDvYaXYkgY+n5ZbnrsBRHLANavoF7mcR
kxJXf4Eelw1fhgGYGd8nfWtBO+Mkl7nsGpRVNEBjeiqJLYAcZvbBvDcWvvb24Z/C
ZF73yRhF16HeN5hHetAmW4gSUVO/j2HvYfZ7YnzcpF4FJkrndqrtgOocuYWx6yuF
bqakQA22hhNm7NxD02VRMFrj3ptdHYP7NCE9KXDNIlVN49SlPpKSCt9wYHF2tRbk
IqtkPIYqy+f1RY4wwdjZgJiP1yLBKgzJS/kSr9tx4YokrXwbJWh9Nagd6mVLOkXE
PFznl/V48C+ZxbEsMlhHIE5335n1lEZxUhbHNcXHEn+fQmeX9udn/h75vVom6Lxd
fQWGmZqjBwWXPhjWUb3oS/V75bDDWxlHkUX2sgmgECRf15BqAnafPwdcvdkif/J1
LOd0zncrTe3NXvEYwFywg4SJcDth4ziMb+UJhIrJWdMwj6Z7qnkO9cjyr4eZ9dAN
TDhK06NRrLLKaKs9XghXZIF3+RrJcRQ/Ug/wuhU4bNq2zCxOgZO1XWaS2azlDrtu
d7oZs0oHCTIr1+dkLQ5Og4bt53E+5yN4tp3KnYTBCbSilUkj/INw4gKIoN6HrjPk
S/AAS3dGbL3WDhgHTXVhTN3CiaIy4f/bcEZogL39sr3aoC90AvLWNA8lVsVB2B/M
Dm2PZXDZqxEp9aqV6/31Y6H4n/ZLWLzZXVcER1AR+GtuZ91lltzRd2rE1rK4evUs
5E/cX6l5/Eedimn1uKUKebKu9ET7ZzU9YPr4DykZ0z6QraVCgxTbhT/a32dbf1r4
graTtEjI8DR/q4RnVzbSFd8/Sjynl1VvIFO1Rn6jXL4AloG1G+NEc7KtPEtPgw/d
PAVxQ7VRhmq/5rQdbx9fJCek1HfA9Ej0ITEmC4idwkQ1/+gnzyPaHYiN+pA1ML5y
OAMIF3u6KIJa4WZpg1g5rDIQHpgIdLqw2veZGYIUxJmjmrnqPZaEkPLQJSsnJBKS
ADe9eeZVw/Yml4x5vnJjXoTXCIEFp7N0mrajxs8VVDRk9Ja49dtcIAaBa7pN2Lhq
jUMr7PvQ9VWlCDQK+aXTUw6zlqefe0JUBw9l1Fen4lLJrcyRjfwDapxYXgEgDMGd
ITHpH5B+yOaWr/ws0TncyAz52F1MGUuMaV/MAhQZm4XmIAD2B8BquQU9/q5mlW0s
VTkXE+w28p/EzCeOgyVy8GNneCMnRkgDOLrGrVLtFfY34ReiKLpZLXuAgXc45FHD
AS66DXBRBh+9Fwbso997D8P/tBHCE2XsCC7xyPhsoaNkLTJgivvVPTS8VDtE1Dno
TKY+9OKmxoKf+xWtLem/aGvmuwvRoNCcuFmJx5K9t33bRm9ZuSK4mOxXHdfoGg9v
0Ap/P3hBjd/K/R2YNU908Ih8lTM+WdQy8h+8MJEe7O8FvFWu8BHLrjfrxxKqiotB
G1Ae/w3UU3c6IDs75dvfTFpQ6IkqX4mOfni7tAaauDG/cmRshJsOKkIre5fEK/vs
YzhtqQvLD2+4HHJnVhHgEd6NA9jbR6rIUyMTzhs4CI2jgzOFaQDe4hkdh/ObIVSA
/YnhjlL5yd5dE5rHl2nx3wEwR6cw8SykOY1fqJoIB4poR1rFZcwylyoNJqqA71bK
x7IrOKQtGnCCkU7wTw+JIatzThO/2mV7JwV7vIAb0btJzG4fzZHmr8bCJLvjxxTD
6zBhEWraUVN0d0FoAbuP9Mpq9E7tv9eBCQ+Cnk4IF/n2/juGQUE8Ulw0EHRK1Wnh
ePLwRPnwcVCjEj2vpcMi9zSarjUW5y3yupDbSLsWkly+y4TA3khjDiVqD8h/qqnp
cJhvSq8w4RiJxAOogRwQjkSUwyNzFcBs7unoHLwKrjqU7XwoTS4VqUowA8qPBZFp
tP/uP27kQDC5WD+aRfNeqnNpNTXBaAIqgmvjgRNr6gy1einIXrzkCLYJemtjRsdy
0upaQTI263t8Q+ynLk4iCIau/oZVl7mS0hgDcNtehPEscnwqHiwurq7cL/BoBnKo
qdx5gXt3NmNuMb/Z/WPbKIdDeZHYn9M87wlOR7DtaMUXiW1QqsEE5Jdrz6cRtKhs
hV9gfiGSiBO0GIJ7bynVDXi8PlW93j+rvx23nBDN4qaIIzlTSh16vWe5nmA7jiAv
0p0vxk0rcVnNkXVvJa7erQlbtrY2eCQOPE4DT53t85mom9/4DDvk8COjuVgD9Vwl
KMm30mr6p5lRUL53qtFit0+2uuz5sUp5LrZi3Yc8O3YYosCElR5rPHD4yPmQrJ7t
x6miKBsfT7AW5hjRmnBjhxeoV7Dj1NUNkLu4pig+/HwMZabQhoIfRhW49ASWc7OT
vDICN1Wvt5iXd6EUGDh8XQx3ML4ydTdJkD9NzxWR2potyT7a57LUFI579rLrLvvT
fVAIvzX9S0kQOIx8jtg9hVwCJCfQlU3x4I4EVvdK8LRgbdkkrxc+KMseKyCHNRo+
wObEMRPKxZ5e7zAsdL3dvvuRljtmAhRjBjn4QJPE7aEQC1NKOG7lL+cqOsJGIs4G
wzj7KcM6ubUTSc1HUYREhUyxSHFaejljQvawJr/P2H+w7oO6+u7zmQeJxXDTV0UY
6FphoxinTXtTXdX5obcbB2Tuf0/mjEI0+5RDNJMmTD+qo4SG2pZQeeMae10ASdop
2v9Dngm1IOwC+l62Ta3E3SpD1BFp3tSaON1OPc5v7zzkxaAFWQuWtiaG/Lw3fSKM
2hnZi/z2MbPriOdLGc8g8HDEitxfRVNMjb+wasn87QhE9sLs52sR7CmqdUw7nWnV
z1FpynBK9os49jBl+HNUER9WElcLqe6SoGcWOqM9fNsXZcAifMd39NGPfPSOx5He
27pEq+xqXUIPTXrRpNfnNE3bpCeQcvYRxAvzDZucgc3VLRLKIwCgTfnrbMfvOYFj
HSL9Cib1ycQboxn9P6s1XwXPma6HGbcHO29UyeZ+hGMmE/B7+6No9XnzH3L1vC+Y
M0h9KkcHQuVcw1AuWk7DX5/6+Z3Ey/4PqwPWFT02oWYUcLbYiHQbZaHbD3ddZDrF
X6Xtj7GI67TLmSi9/76lyHgQsaJP5PcLIyfMowQBSQbnQnZtBLHt1Xloo2R6N0JD
U0szUF3DnOVLH1MGZPOnb+Q8BvbTiqUQP+toQQKLHHcOd4zS7TX7pEp6mWwdpv2W
YVBwRKtLm8CtkW94ArQG/xshBB6WdCEhB654UMjrVjFmakl9h8nKrX9LROUaOgj7
7vGFuTNouewZbZGn0c3NzAhCFJ1DagHeQZD4l4w+MoVUDuytQ/92RHEJFf6x2VOj
OdYE3LIHJ86vRMsC/bMYtUXJILFsOHc4wgXdyOUguDXgjonc+fBnCj0m1u/VCVFd
Cy5wgL9S9FaZFlLSbuJYxxJjICx15JVXT7N55rE3/doMfKx4lU4eFF7M6XiV03/3
gBXBokNukrfaBBv/SZvVJPDL9h9kj8G4hnmNxdRTpwq13mQMbosWnfH+jJBEja9H
R3VmGlKCSr5efFTe+Q/xbs6fDEzCuau4kcIlcYlmIIBkUfajquF2rJU/ZwVqNk4n
c9pzLJ7tNiAw9JOOafU3jeJ/G3XpgctKHPFdO3STDDxjZROvjA+IK5xNBZ4aRXdH
nZX482g1KEfOMZCmeP/GAdb+5CLsjCOSnRk8cBivhUlN1UXY8jLMCpUbKKuVShjT
brsFRhbA9lftX2f3Yl8VbrdB1onfMY2aYIMaQypo0Cch1A7pUtNZ6kdzPs+Mkazt
NRRD2yybu99Ab2jZ+75uRVMVwYBz1sr3fiW0FB7IB6d3YSHcQsyajHigM+18uvSW
UkaYMMuY3j10hS85kZbzEDMuSTQU7MTYc8T8D2SYWV/A7CoRihGp8oGym4HkyU2r
n/zmmPlmlbII52otsnzA5R8JfGzigreSx582AmHfxTonFx7vu874cSJQisueVI31
w5iMrGSi103usD8Y4oy9X+j2elID67KKo8ylZQH15u6664wKPhxCP9X5Q7dwvZyy
/S++eNnzLPR9pWLGsnZ3mW8R3juzuTJxUiah+ZQ8Jjk9eqsOGHjj7ay6jjikvcxw
RmgCdIFXyEzRJZaLfncehCHJZLywPU/YytKAvuSY45hUfmAZaFptKqkLuzniFUez
o9D/MZP1RsCY/Qqva7vRUiVTQ8kZCc8taQHh5n2B/i1UUX5wvHcK878ACMsDQkHs
P0kN/sskSQC1iIBXpK7gSwVmGx9x/sGbN1GvV94+Bugi/ds+RZcqqCo9n2DqJ06O
SvRMvT+lXcfw2r7GpjpeJJEYlYVAKyVqV2ExUdK6nEway3qyD/dnkPJFTttb58oY
JdCdNePS1Tw91yaJmM4lTqLDaZzDIJimIGsb9IeHRJ8l+ExpTBi0gdgkkYQr92jZ
AB1kZue7JEo9WvpqPH1hqz1wt2Rr3lzAabXXgDDredFR2K9p3QvKT6Ucm7TznM7G
uCBDDxmfXY72loPtq+8FFoV6BCGGIw3RSjepKGatfK5rRZ4iViuTpEwyNOF0HFvQ
jZhVz9py982iQsaSicdLqFe3yLXSODO5O+keLoarAZwkjb+VpuZyVrm9pl2mDbkj
GIQczYLi2nxtJYkj6WwLn1SGX0IF79XmF88j8Krxzq7pL/WcNWN+7L6x24p/brdT
6JXjcb2L3B0w7tVsiE8JLQfdDF02MxErmRuDtbsgsyI1S/kcDptpGLB5vPW7RjKx
HL6mrtnzf3zZ06hl5zw5qHjFtCDPMqxGXa5KQ2/7PWvhlezCGRZtfNPV8Zrn676T
sYHf/Tk82DjZ16esYI2xafnCspplOdxsO4nchGpiZlXV68IMGRNW80N5UmLJ2Yof
2eyXbniCK4QeSF35aph90N1UiRwpssmia7sB2iPEsXYlSINXQGmZrP9KRDc/gJv5
fvHGgU16dfmNizzKzBzoqh9gVwc+9lieSfloYNQCE1AY7asBEm+2VJPyqzSBnrQO
MZJst+KnK5HeaUGQRcZLeWb4YMVesoAc6wyvletbNYyNGW5AryEwpTHh9CfBBXZS
/g/w7in1LCRw7u3lcADl1OxNUKvNNx9n95u3fXzyNPLV/3XztmHHIWobzUN9wyHV
D9Q1ciRpwSTsJSzdHfMp90sHzt5fBWNIeP+twQ+snvOLkBGymW4/OAyJ+P/N2ip1
stFSiHzhi0rgGRVZhmkm0UpjfIl3GQJQeIj49lQi9gaRMLwxg3clzQYI4qJ8eMzB
Aj0DNxq3+ljD12n/GkOrbBQNLE6hSsFRrUMxGtfHPBrzA0kl8ZJt2i4bI9/hfEd+
P7Iq0RmpW8GnVnEDRsUBFbOx8HhVjxlV5M68LABtY1yuLAA95zi9PezVkVWLp/vB
9Y1H/qAstM7s6UshiI5XK+Ycfwqup0kiDhi04ak2pEpLJ5Vks90ONBMFA4IfRs4u
AspYG3FVpl51zEdtM1peR8U15RflQnUVrFxU2dJ8ovNUX1zPL1LC6OhIFwq8ZsKj
g6R5KpD7BfOrECFwVKiMrubtfLVe2JDN/0leTtL52iG+/VMzpVnjZwYsGU1Vvida
hHuZoN6kSjbkt1TLuOF+Zlv5ogosYHsK+6FbxVlYFbr6AN9jI9a3j6+ZxwanoXqJ
KqYvaldQmbuD+g4RNHQ89DaxKj1fBV0TXTbduAh4gZHtF6pWjLEa2hDZ56mlbiFJ
bKQ7GSZ8zi/DtWpqjIp0ML98Y6fh6jz0664gv1ouudHAlf8GGV9NJugrCd5VzQ+p
U/rPxlwqgZmsf5MeHyRdCuGw5Jxgo3VIPPLAJTp2cdKaSvFVCsMhrOKOyVk6c31o
sqOYSzUs6xykGCQnLb+Ym3E2HNRDx+5Pd3MDV0uS+I/AMv7ZSpbCpcIz7NVaoyqU
j+eIOOfK+J7Os67EWY3DqM+mJVhEU/cHwiEosSad6c5iMw2g8ougDVsKbu6r4HI4
6rF0ovoEJFByjbFc+xsl0wDgw0qAElhmG4Fdrt8BH0uREbe19hiCIdQrf77qIjG8
J0kRrXov6LiM9kZk716IN2jAzHbgUfxeNtf6TjTClhaOhFEoDxG0Xs2ler/JALpk
z7V68f/JVLFf99MDmP9kLGdnFxkDYI+H9JFOOyhytgmjgSsLUDlljiNSFCc1v/PO
Ix+saqb5RR79YlENP7amaFeCvnWQAZ69Gqfr6nTPWqOcnxIojX3ssJO4MS5b31CG
q70UVb8js6qOqvtBxUyB6edsr2UULBxJorX7KAbm50y4sbBmp0ZWuRO39newgAb5
XACiIPT/4YI9OvQGmcJMnhRAQhdnTbcUL7guHxr+NAYxW8CgsLWGs6PAz4mlrNk+
78KvM2Fc1II7n0JIpSgl5m9xEztdZrGt/sFr3Pe6BjOiaD9MMFL0gKuiQlQsjN50
kYMcGSqyERcN0RVB9+mfzRIAp4AbgSodf+InM8OIczqPui1jnKM/g07Q58BYG6pt
b/0Nh+SatB968dDyLnPlwYWe6mbmNcpUpWYbBDTEtT/sofyfH2w5epcDPlMLjJ3J
zoWI0ofXb65JByR/SGnm20c6xsoE0G0MWDXPkp5KjJEFh4lPf618VqxHc5WCf9v0
/LY9s5nTC7QM7NNQ2qQkUTmaKFQI9x2TW7HrsvytNhMVhkeO2B6il1GqB9KXj9i3
RnuJbwNHBrMUv2ZSAEYbXlRwCwqVCJQtL1+24aHVMMyH3gU4pwPHgMVPxGCHniGN
CjLbkTQjrqckUOH5i+R/pXhtpQl3pY3RHj2ez4ptVWU79fZacCTYqw5GtrCnnVXt
C/LwW95Y7du7O98gB/ir7fwEH7pDl4EbmJGPTPerSAnXDjKGfXwcVn6CxqYWEiGW
B87sLYo2MTVAUtprsIUBGu7S3gNV+w7yHpIpVbx6m675w9tJLSab2W79Ot/6b0MF
FeVa9tntnhbirT5g7d5OaUbJ9m3fq6ujtwY+Sj/+FcN5kPKGEH6KuOQalGg+9Uaa
g/8qSeRbo952Ee+QucnzGriDpmE/ye7vHSlS1kDnSzl6hRErLgtBq7M+j5W1ipTa
/mGnTVuvLSlBdDiw3BcGj/ZiQPj0scJN16g/hlNfDwatA8hk1cx/HPbR0AccDWul
beOvISt3WIfKXHv9thvLqAh4wo7J9IRW6DMYM70AcCo/2S+gg8PK5H8MaKHjMlyo
ZWn8DSw71A2HtPhIXUm20Nxb5hIPQQdIkAxb5uJa51vBv8GzLE3FznI3iHfu90VH
Rqk5eu96TLfCNKBHRA/mtqmLKuyHktZJjhbvEnu4fLUZwkDOot8CvVTE6su9z3+D
1qvSBh1MiaJcoDmvUHJBMVN64VwZ+D0N7R5BDla7m/ECt2tBxdXIJhX1zigjO6GZ
2tUy+oEiOZJz+7X7BQkEQ+hSNAm9ZGfWQVSQTKcAiB00wGDoGCdeR+tFi8vefJaR
HBXyEEGGBHNiHJBe5ZMtlC9ZGVh+QvqI0uj9+CszI2fdfyzYzhxOwX7NopS8jF98
uHJE/B5ZGQXDf2BlXObKrmvMhpxGqe1RhwRYiUUUGxzMN5MMN8KC8I8QN0R8Bju9
C8Y/G4MjRosgyt4+l2MfMdne5eQIF+h6PF2acyeutK0uE6QbLKW+FN4sTHh63q7U
0+nGHlUsZ5u5CImCgjn/a4++fi0Wl9Gk9xxaPsmaT1DL5AJig271ELktOAK05FPb
jnYMkqfDciBKOlKQMwpiYvewIv/QNDf+VRsanrPHvPfRI9cyD0hHOrXZgiF09NyO
Gv/qoGwmO9fAiTi1d314b609eUH9454C7aQcHaki0a8IEUmN1Wptm3mexUIWxAHA
VOlhb8/yUIvQUQYo43n+ojv2XmpSoPidbAEwm9thsJgEC1B0ZXxFI1Qc2czpAfsl
c0PPdZmnwCNg19eK0TBpI4EHUZuMZJA9sLZSu/cdm4RPgUs+I/6LaxLUTomeLGTq
FzWI8iTxO+D15A38wfchQpZdjaqI5ipJVf3yd6F3HXgT4/cip7XpNA9cz6IM3zz3
YkBGc0/DVNyZvXydUms+SVb3YQFaMVzZvINaceuiMegr6qs8FMxLrQGXz4g1LV9+
aWPZb1kJMjpaQRS7BxVZFRcBf35buqrPg2vSH3q2C7y/gNZ043ids9MgDxxwMysg
UVWzk+4w4TbwPyBw0ITYayRlivpAjphn82jo/Ik2/c5wc7lu5xkIyYFTw7pWJiB4
/zuuST3kEB15HEoYsxn9U47v3qkRvJK4R//yxI+Q6+V+ohAR16OhWvVtGUGfnb1E
lO+9B+zVeFbg8vzIClVfU+8KpOtjXg4SYYh/AzadAVbQfFSI4gpddDYdlP3mTfCP
6ElmHQv85AMHXp9hGTPun35/dnRr0eD4PzvEbzKiIftN/Jzjy/h86NG7RKECRuzl
KLEQXFd9lylV9CzSpusdukfcuD8P/ZV4aWk8ezD5NNLO+ZkaiFw386jj8tq5gNr4
1I84XDuza2O7CyyA0N69HlqmghubTMrMoOVb36DfSyI4jT5lWAYodEo+ebHCA9v7
VCnnJb7PAAfz6t/BTDKYLM9ZY+Z2qIFdbCfWbfgPp6P3/t2zQtDdkS1+UrXPEsZT
qPjmnuVeM+sYZI7C6LUcM/SfCrsxQoTFT4p3jnHdE2k+D2KqHciQ0nhiO3UvQ9Bv
E4L9YQUSNvibGXJaoJtLYkdgGCkwumVq5tx8936/BNRLPWSADlCesin80cs8wBtY
gyHwvNVd8OZI+d8UI05ghRYzVL6IzLCTAkjnBFrk4AGx4aa8IUAmr5/TnhKYFFnQ
qYt9XJYFwMhiWMsFImUafS9dBD4At3bl8pa1kSFNJF5R6KkiFl/sS0BH0tWIF+fN
qFpwxt8U6E6ynHCbvAHJtW2Kz/UZ5T3fc5lIGTCcdR8Pv/njGtYrQOrL3hflZHV/
ptU6HI9ISbebD86rH4ulndBM8xGmGd38rHJrsqzsfjf31T5AaWeI1ssr6WU0t3rl
an/wxO/qarO+lnMqeG0oxePxk6LKqN2WAloqTG8wZXTf4RH0w+qdJH14D/OYgWYf
2tzJqHgiS1UGoqxbt/ruDX22iypf2UANVFutdCQwbKabDz0AqUwokoM7G/4I0847
jE9pzRoNAZI8ANWGLRPcYMtcW5t9p4mr/vj5v4jkcJyOwvDxLOMFpjNKx+Pqm6Wz
ex7ISAo/yIqJxBZc3oK0/YiwabbyhzvYdHf1TEg9lHAWZgX2thwiErVWEUAoOXLa
eBhTzlvbOviTrG9WLX/hQi9fYs6jOtXUxJHZXwVxFOKBDpDQ4I9keuzCoHyfi3zi
Kp52EprVBVLXHvivl0DYT0H5yYnKc3i14DQWP6kMaAODxJTYF8XfQfwW7v0kYXnw
Vq/2hTO2YcgfeApAF+RUZQ0GmCfkoCw0/w/M56OYxa+tHWN4m7K34zlRPFjpDs4h
f593NLEl/1sNE3BkQt66YEIF6sUqVYeK8lifOsdiiyKfrVjBZxsYDGiH70KGFohR
vRJlAjqWP/wdRdSBqj43ikAAn4PxsNsdC+P2/wRVmjNqb7/U4QPzHmFt2jUt4OFA
ehEdfjjsMHJqUfX6vvNtPkh3VLFh7AVPY/RWn6uC39wl9pq7ulQAJ+yHCbhoFBx4
DZyoOGD2oSwS6A5eZC5pmdtaJlv6LgJ4SRneBRKNTagCKJEgQvLPZYta6s1b948l
mTK7Igb1JpLgM/CLUe2hDCEnoh4tTNEY9SDHfuFyQnhHdbYwivHZp9q9RU87lQXC
17pmoPs4ZMM6DI/cFxD0dkJt2qK2JOg9cVtZ6dD9QGF4w1SFrBbFvDvEanap7WVt
4+SMliW1UkTguV4RbnxFLIZOQgBjbbvm5ydeA4o5VPHLk9yTrbL8kh2rAvnq+g0E
CHXWRsI5RvXOWJh5hEiRBG4RIJUaYSl4a0OJ738dPUw/GPAaX44spXH/pFB1gyTo
nb2P2Q+taATZpk5//MsFxo9NnVnGjx7LptbJxEEtfRW+T9aLI343pm+Wa3s9t+wm
nX+4IqOTr/4vxnVeLns46FoYdme1mNc8fL+ePL3l53dkzYQFk8xGsYPV4IjWy2dv
iM8neKnbaDIA8mAeTH0JBT8kKAXwzEBHv2vepiNtV+flej5v0FNJ4+xAuCLlW9M8
LA1oT6q+WBCq+wffuiOXAOoVN6Ow6eWPDPfCsj6bIcNejjsyn44cDLkYq98eXyfX
cO7mCnzyobvmr+4XVrbx5q99XK9xdFehivoh+vvTaNaSl8W9gtcNPg+FEiDQIOac
lv8KqhVgKFmjUNU158c2EuHGAAGzDE1KHKDfgRXLt0UCf1Xw5xIcxzDvsEjm9u9c
QAMBPtpaJtMS5rrJgVnvuneNVS8VHMvvwbFpew1vkpKmDYCr1Wh68a1B6qbHC0W1
wMiDipUzuwINeOL22teNq4jl39l60XWyFvvb+O3iNGMvx/S2INgp9X4KOCA9E+qo
RGu/onZF3hOec089P75rY5wug2KLKE1ttg+812Bp9NVckxyZvQxk7d8qKd3R9bfg
Yo9S3iNBt71d5Wz7hg5Ph6aMY2+D/FpnyZWMlIgfo4TRLK0AKcdb9WS0GIr+EMK9
ioB2nVOL5ERF9hlOFhEuoQSn9WNPaWMmcmfi9Ris06+dmlPFVxCZq9Wij4/jlcy+
FnGsqOyjX4B4TnOskR/dmyoF4N6aoxSqE2D6NSTU01tQpaGvwo5F90JfD/3v4JmS
JJDrDj8TPZXmi6yYrukm3hfK0G6c9b+xJWGmoUxJr691y1s++cjxMhK9qNpcb+R1
brhyKflGYfOavL252skK6OxRY03zq9/s4JTMlKu3S1V8qN7pioxo10Gp8j97aLuh
nMMnUi77ghHkH7fGPdAOzk+u7P1SHQrdWV66BtCUYPVnn1vMdFgcoQpIRtDcZLPV
SZarspUm24zCicbM4VZl6/EDQSyMKEhlsT3LiRKfiAzDY2zQFlbsY7GAzuLSaoXm
OoE2BrR4xd39h2obEe3MP2RUfiVufyGWn5rJpS5+vazmLPylzZ9i7c2uQkIhYbWd
ONJXzvGgnAjBF8q4H7FApy9yt3KU+TKu7c1RkYyOuhNDwEjsU8tJ/TNCsXLONIrs
ifj8nboF8xc1WI7O4dakxV8mzwgl6Jlxpc5vjNJdCt1JfUx0P2XtYq2j3fKryOVO
p3+e1dlou6F9Wl7dvH6PgmltrbdJK94/469oJTgBQSxCbbNr0L2phvPfDfVsikpI
irzC15rtyPakav4mRLcCja2/vZ5ED03JugYoyz4hZlLkOESjKyBt4y80sL5d3Jde
lPZPOp4bktXJkicQiqCUotZVEcszv1WBU9BCANX1uxvJMras45is/xxZDX3Z3M0R
G74rLojPyoG850SaobaPi1L2ObQk8XgELwhn98L99LHF29/qVrR10ayFL9zpPnmp
LeBlmBldqETXe5/1DziLv+NdP6UUQfcG78e/1IRmcxv15z+MFxpqd77qtzkAdHow
p6h5Nra/Qqmd7i3WNfCjcrcJGN4jXkMmVJGjM+HrXGDTNxFf9dyCaI5X0IvPxtUL
1yWfskrqqNeDOpIAdfb/zLTR3tf5Fosl+chzQp1JCm8MEJURxYR8U7Zzja2TPJlu
R28JOo6fWOizQxY/eawy5tt1jNNZT9Cn0WJSNF0SLPmOKzBBgN9gDM0kd9FhuCvO
vNSg1gxDCQbrT44ZtBeK8oDvoLZ4QqUssFejXK9b2uOKolAuVt2tmQz4L9s6PNvG
/2Nw9lNzVEXsAxpYl8F7Z7leJQ6vnOr+QLjXpsqtjxY+THC/8Cw2JwqDNONWWa69
9rUX7/TCmtRLlqFHjNW1PBObifBi7I0l298iJYYNdFWXgBzomyQs84PKiVNwdJML
/hSVDXvRSwnpk7YkBNypqHrPJGkcVpV28gr6owz0Gh/NYTaftL06FPCHI6UqNggv
JXKArQWaBpQ0LRS4uoTLMn2I5zdZsHBw5SS8B4oWIGgYuZxkwemNh0LaQkpppm5b
CZmS4hGDo4DyD61brDtw7DsgSgrTxK9y1oXRibXPVngmjafGruU728uAaoLDdqDI
QKFg1B8vUb1ZfrTde9S90+EaQV7vV42dTR4mbUifHy2P+qRQiCXakzax3Im7Ucr1
Myj7/oBcMfFluw51zej4LOoNngizto7b+WfRlskTEHitm0Bi6hTmj5RLbaPxR6/w
DoiphlISfIkB1O+NSF2KXj7Buq4t2fnqSfqldZdpX2PkQ5umxBEuLP8qxdv/GL/w
7244TBcX+uAhhRtErRjdkRjKXHXaXcoyxL9YGXvdyOy2jwV8q6sTw17PiF02jbJ9
Yry0YBZqYcboKfuhWQEzkRh6v10mW4I0b+sD71BpvA/iScCOjT13heuWein9EfwM
2QClOcIP6zhJmXaV4BtD8qTqIeXAifcvJ4E0LBgfG7ajYOzLYx5XwH03a9o8kTKT
IplS3d1EYi3W5jDXqO9/Pzqmc19lGu0kX1Opgbwq21+/w1Kq3vU7lX6vARoqr8QV
ddb8otR8d/Jmfri9qwu/LLpgzDbXMLymIe3wcZq9h0cNYJd/DvqwpuH87ei1Cs06
AAh/Z9lRM9MSmq9tV+ZRkhzQpPDZUhuI2abH10gmIjhvGSR5xbdrmY+8Gw7XyGFa
c1WLld2zw/pvk2jTpptPf5ZMsMQaaCyg30eTfJnZ23+mNmdRXXC6JFypUrxNrZAn
AJDdWHcxcFOEoESw3zwwxwVGVW9CTlxPXYZe3Fbz8myy+TqMyEb8S5xl289mvgHK
4vjx4S7h04R14U7f2751kMxj7KFwyKpZbY7NboN27G69qLasTyhxEnP+yKlvnbTl
dHbXCl0kC31ecXPcbnmndLnQqSSW3uy5VmglJlNGVAYJO6UN2gBeiTGW5PbcAI5J
sOmwuM7lIQKl074ZzyzDw6FHm0r0MqrAmSuFm3A3ywIzFGxzKTLhGhxSEtiEJMqg
B6URND2DMkTck1lhNUL+0bUsHFtbstGbZs9plmMIZOgpgQXjCVYZ6qWODA/zfrjF
9Mj9GKEkgJWiqwFac1W53CCMg62nGLBajZ2rT4HAKgvJf1zotoGloYG7nxc0ND6C
vGpTAxigi1blPahNwUtsigd8UxgQj0TJADtgXu6QIJxoQchvt4PlC/G5/zMxx8/d
6j0QBYfMNQeREIjCY+dmqlRCp1vFm5ICQBNtqb4T/kT+nmMoqI0VkLwC3A17ZecL
qUOLrsgOB56khbUzqqu2EyiElAA+sw7BuROLm1G3J9Jc9CR635SARZnVgxf2Fei9
zSTzC7gpkOXw/rDFB1YxAbG4plNSLzmViYRFDJPz/k5txarm56Qhf1Eus8+7ecj7
YwCDxmfQiTGlXPR+ZPC2KZrgbk8BCuIQrzKYpTH0s3FHl0cjx3OUxv3vzZu0d/Bj
UlumZp2kQATQopTbaJQkBKrCOlP6ztvtdxrHHRo/ach8GtnqPFi+VtJX+c3JN2El
KSjIr70HbMMJpa8D5DpO61DaVlyHOZEgYD3oyrBO5uhIb9rUCxPXzOxHMIxalfQT
FOTpNk/SEqt018OSUuix8FbX0SdzPXIRVoPd5E/V7urP6TfxowsiRlkmavaGnvK3
KRusJ5uPw0DhTQgFAVvZqD/WPvvUpKkMxHEl/Mid9ArqfLqd0BHCHgCERJatpZNs
ySA0y0sXvqYyoH5nRQ3STM0cFDGh/Sy0h3/0SlN/ihwpYVFuy0JYsClugEHOpIGV
pfWPqoqLkXPMT+QKBaPVznFQtPnBaa3bJWqAb4IKMY6BFatzbipzr7bLFMtl50NK
uYw92ISPA6hrSCT4w2pGGD38JAHMkZOm72uKsfKMYpPV4+ey9rfvo3OzVtRtGoZj
FfqWxfExe+cl2md3MtqcX8Apipy2WtxMskpZQ2SZ6J0jA6Dp0vSTDUfLqLvn+WGq
QvtAwL62TnikYngh0DKM2yzpHY57uZ71SHcewl83gJeEEZgw57BPMQ4/JQCrhwVO
50Yj0rAkInKuDddQwdtGdAGQluVYe5xK8/Lq+y5FNKi5cw97aWkbXACwJGdjMEWV
PbN7I67KplRQcYHSIaBdxscN2N7QOAqlzo3YZuUsKaI5hAPjdso0MCv2MouLANWr
wUG0i8hC0RD+STzbcGJbm8QYQvv8YNKpeCRIVvQbThpO8Ld2cVkl44+xAZu366bt
embaxdm0Zznyf/t3q6MEyf4Ko5/znqQVNXP/0/hz+bjqVwVXpsghNpQ6T9DNCITZ
lniGG/GvnHUUHxEcLOi/t5pS0qx5/Zftz81O/veqEpzAn5b9DrIyZ4YAfi2bKHZ5
U1w69+SGi34Es6tAPFLv0nsBFN0iwcs9k66QwTFqIF+rRebZYtch6w4tSqNk+6p8
12GvIpgTHsu5ajwfUU5K0fMeymtnwBhjrqD+1RBGvJhGpawQLsQtdFBzLUKy0EHH
IcJyHbeYHg6IquaOGfM7Th/6NITHZ/l7LhWjbhnP4hRITTJL8Tgm9pe4GVSRVaBe
B0s1c2prIkouXF1dlcFCc7QoNfVcs+xDBJpEUCUFDE/Aw/dm/VLT7ZmKuWwcG0SG
g0wrEgnmTfQML7Y4JtDO3X6xXm1er8vrHihQKJkwMDaEoq2m86sh50nZWBu6zyAV
Crmi9NoXMys/MWO0Z/rIVyhGI8vTyr9vKGJlxOyTUqYtlCNEiWUP2v8UKtXYnUA1
iS7N26zEDFokdJIr7c0vc+2uv6n7TIftUzU6qT5gpr1T64wgwI0tM072lrkX/O8d
rBrAwKxsAtrr7GMBlKTfrb/W+voK2LEZFdNo9/6ZwLzTBiAhWesGAO6PEnYmRgPY
y8vW5R+6wb65MRs3D0Yd44SR1qhuUTobN2VlBSpDsa2sKNi9NZ9Z16PZqzqiQVPm
Noj4WPGc+9cPOipBw5Kc/GcxNqKf94avLntkgD1TavXO9W29WJNCk3DDWgVfrsG2
30RKazD7ZDAiKqKt7VuDwzZzM5jfrMPtAgYjmlO+yNNeucfX/01JuP8y8ae44WC/
MT85APIqg9QToT0/fXrJwofYldHUPiofsQsk0+Y6UIXwJEBcYh6Lr7TIjHuDLI2U
Nmj6RnFlV4GQa+pP46QHQHfoJBz6ACa3+uOoLcBLPEH8KyqLqrUldsbQl6BtYY5W
Ms2rZ8QfvZrn65NrMz/syDNm23zEtbx4ZIMnCuSdLakq/K4GmBiBAeuvlgkiOqIg
mMmo422dxCN6XCvTmFV2gxvLTnEUqTVHOHzxwUN7X9A/gjc0Ud4nqEP9tTqSXtdz
b/mJ3kSqbPg6PCgiyJyKr60tzIXwNH0ToiGTiH1PP0M3uU9UleOlFXEl1SpeeoiM
sj/xSIGehkVImcNeloq0WHraK6ZOUj+boi4YQCwgv7YP+OdDwKMIyAc0Wz6d1XW6
g7Th4hKIRONSN+2ILZLomV2hcvFiD2PEKZQurrNt+piSJSJVmhXx1rWUGMvePtT7
t76e2VxzK3Q8PI4502E6yniai2XDetMs+udMdmFqgbuxqWcf9B4skpTQTqyFnQ0M
iX4v0lQeb4Q+3UgXAzL23xBIi1Q9BFSeVjzBYa0qbiDr8EsLGJfr8/MK4Zv0epy0
cE6p10pJpgyAFMK+VXz4UXSj4Bol4VDJn8bVjS3c9uqz8UXvMGsdSNdxOGkE4Ovm
1apk0aNRdDsnrqm2UO4clkxnGNVE0ZwcgpH0gFKdWBUWk0XxOfnE9QmkS13kcSW8
GYSBMsifAS8Yt1O9vZMwuC9VPFXkxX2ZfRm61IG/xZjFzY59Fa+LRN3QZmTjhAk6
YuLAHpv9wdtA7KDIc5xl+Ca5b7kLKOkKMf09sv+QIfoM7vc4nM+0rwvl0v1bQVa9
SODR3jIEj0ITFHTT8Jy/ICMQVHmUlNMxPs2lA6RNdw9gL9FzRGYtKEiifQnR0+as
tCJ4PivPzfB5lZQthel7YJS70AbL5ckv5EIKSyKmy2puCbOIfLz//xEbSQRSaDBP
nb26XRiQpZWzhoJeJYUFLJUQIFqajsyCfiQREmTVVJDbIwclPklIqEL73mGTXWax
oXWiK82hJEycG07OQHxG7a/6Z0PCLTslmryHNqta6mhkzmMHaWE6PxnF9HQ1u69V
UBMkcwvsPDX82CtLU6RhnYttuKJxgS6eZoKCgzljKJ1QqQQq5p2z0/KXLvGWIyDG
0+nVOJkUo73AsgiA9BMW7e4+9+szBXoXkca1cWuiELyY/+HC1utrGwcfAPSroQ1I
1KVfbvIE+D9xFbTEyYgOUUNxtSJ9bN1aBOb71EbwRxPbTAS252d/hyM56KQeYBRM
I0p+0rxJRPn0P1C4rW2OVOx+WjNHZJvlquAkbm31rbMS5GmCle6zim78Imd9Lz3F
DwukIpnshjvaLK/feXb8kWLRbXbOMYA0KFJWFw2/SV+mQdsF1xm1es2pgRTvcjo6
9oJrgTvDuXZLJPgLyzBm7kH0inmljeQLp19rfRYowE51uiqQswjU507Ob+GHtj8A
bokh+AF2v3LjYEO0bDNo7eMwuBRTr8r7Cq3o4Xzztptg8gGIhhnqMwzSJQjEa6eO
p7s37QbKeJxeP+gqajV1SIayvDG+BCCexNLarPgLc41Iwg3ybKWmBX6yyJWMXHkY
xrdBLs3hup8Kmm/8Mil538Hu80jfiARY+XVOxUuLKqbq+eeT+kNIXigb1Iku9M81
eF251qaRuhR9z1RpVFVGwSIyJI2DCF/ECiLWotUwidiVhhxmJbRTXn3dfNAKvqvx
NkVTHQX9KbgE9WCCNsvistr6vYmEpuKPowIIEyxNtByG8qK9xXjHQzc8SJA2uAdH
5zIMj9WgeG+HzzVomsFNhrM23L7x9oF1B/vjz1amu6FMPomCnPSzs1kc2hbDPqvv
fXlVty09GxmaRd53TLvm67LDVFcUY8dFMBs1AY3Fh3d98gX5msRK8JQXwwHdB+vW
u7AeOybXAy+qx+BCG2hO739estcCw6iAudue1CzV17QF6xPSJOgpfMb4ytTLr4Yh
R94VTR3rRKrfe52+zN6SV6b/uI3QwIsED6ODCVkO0ZjYxjELHAi0RHcFLQHQw3Tl
+CGJRFDgwxqfYc9JnG+oHr8n0Omq9ypj/6try2ax3xs+/CmupJnUediapGosSlbR
GIlb0esRkI05Yqjgxc3hz5VNOLL4HNUOgqFA+7NYqmX7t1bsBCeUp3n0RK4Hq4at
xW2nymPPg390RebpCiNSN5RJHQWys2nYaWelTkNt+Zc8+86RomJPxl7KNve4mj70
KVWSlmhMTgqb48JrjQA1s6emuOZ0YuF+Vrgnv6P1OCQcc53UGpul3Pu/Bvak0U9d
s1ODTPBfT9DepJICzpeg2JedTGnUnQcUwPsKfS/aM9JVRAefJlHsyTNJn/VGX3or
B347UVRargKW49tkq1mG017/+f73VB2Phmx7cT4/G7lF6hdINL86/9FNrbA3bU63
3WJQs1kmArKAxeQSxomKv88A8gJJXFz64irieYptzqzdJHFRQd99VDJ/1vGKwWkI
YPV5Xc7yQK0hf1/sKwmyL8D3TjJVKr72xLuW0VKI0ywVA52jT7MxZgXs3Z2nsPDK
ZrSN0xBaUYVoiq32yiBLICtWTaEJzlS7KHYznAoBkiVRm7vj8w+FetgXprKkyET2
mdu5DN7gFS+rUUFATE/My/z7dOHV3lAR9shYBNsdRcQGYPVHnzdzM5EgoAmhiboA
SWehziiRHlLf9PTDJz45qincPDEjmyISGp7/sCwkQ02bL96sapymK+BrE+/QolyO
vOXz3Oga8eJA27HP+ZdNCaH85S0/dDoz41YoG1376otGQI6Sq1y8i77pBQpO493p
feW8sEnZf3NNl/COu+m7HkZDGThAZEXhb8JBTraixBR2JW99G09mc2CXDP/qNt/H
YoY6IuUgJoNUxoPff8L2V2cA5QMu3n7KJWrQ0dEqa1WSKRoM4wHFdn6rRepygI8S
TZuBTLenKKWME52GXDE6xUnr7vH8owYJinfpJx0vxproxEWd59bwt0itrVpfzH+g
vKfCnWSxEb2L98fF6eRsZ9S4naZmFI6l+QMRcTa/IWczgFWtxJLdphMgcCG5vmHf
di8VT2AhnTPgQWW/y4DkWgUcbduqyct5/jt5h2+Ao2pNDQqIjJ5rBKK+Xw1lGEYk
58oQiXxvPG4HRv0G7yZHSAq3kyvyFvzMTNgaykrWpzcMDdIUlqeVZJz/CXVZ/MI0
PVQRarAxjTLlNbiif/wkFhdgMkkVVMkVplddjboaGN/gb17o7YTgcxCcA90p6lac
ztOei8nzCahbKF4xNYW6Tu9E9XZAESGu1Jq9C37UqlZVF7eWbzsMRLTpLpNlSwp8
ls97OHusjyAvn4TOeAd0yvKynPO2ZwY/j41oSCn+Ox23wNttKEZ3mtZnDsLnks67
hlFmyyKOZ0JZycA+pKLn2ngOZ6hj8bc9aGrwC4Vnc2euyVvCfqDoYgiSZEncTWhy
zbZmBJGxjUkO3r6NvYruQ4AXykm0qVxYPSN9QCQVIxwl5XkkuW3fs3wBsA7w/cTL
4CQHaM6Nu/7pZG1RGobk8Z9jraC2yRLnYPQCBmDa+1O2ag+dGO5q6hOSyBy+C5Be
spaAySTDOJRRQMt0mKxzRDlTWiOniqkS1ZFhqbKjjwHAQTTnkVgvY5osxr9Nk/LZ
q+AFhhOgUoKZ/zcyosdHLhGyDxKVa2oYy9ya4pDm8IK4oG5p6KdDyBs0xX1OAy6n
o1q3xE9L0+LR7EhqT2YjZQu3XbEruwNuWIPvo1QSWADzcijppwfggqTKuXjQrz2x
TXc3BoqBnADN/z1SlJ0KEW5cUBavlv7m5JbOBi4jEeGdsXf4seQf92K0rasrBNOA
bgPdSnEMlMGW0FJlRmZudW/WruVySRcuMTUWYGUySLnjZ6PFJzT9DHyRQGf6xele
wwwWgJNgzlFckcqdIDbWSfGBUTQ+jImXMa85FrhcOBAX7EumQiI0LvjlCbA3hIhv
ouvIBXWweof8L0V8W9bHoFp/6NbyGDVuk34bOrDPaATxdb9T1+6KBTlpKO6H7ljr
ZlyJVcOXDrmyORP1PpwdfnzZIUqEaY8t5dS4H0o+89dnWLtLqwEdbJdAAvRGYfn4
fQctrclNvMYdPMQZ2gVblSH3VkaMu7o9UPIF05AhRcEtkI3fcnXz0uuYhAwMk8LX
vycGO7H2BRW3op/WyxAOpcqs/6bhpLusVLAA3+7nyWk92hElNmBnkhcAui4vJIPn
AxAdupf8oekW22Goma4JVcgwqHwGY3Imf+LlDtRAZQzBO580ELXvzKQP+ByRRjmT
JJc9xbCyNKD5weawvda93Mn6D2F/UJSnc/804wXwoR6LGE4DiV1ICAHiEbu7yd2p
XcaedrbrpgEcpQFsyP+9SO7SYYsP5PXnarvnGHBHWCvUSttykDRPurb3SpPoBdEp
sIdhdmfonXlx8mQCnm3a2Jv7Ajqg1o0uC4qjSBJafu8Dfsp7H+7dvQRYJGffTC9b
mNfzqS5wIjDMlhKQ3EMXtPkDauno139nBA1/KGPVCUoFuX4vXjnFnTV2f9bbwKRe
QAgWikZMpm/3w6mNxgFnMOeiEpVmf9YhqOBWWmgrKMz6g0UW3BvCGZhmwoqa6roK
dkGxJueRDvLuL5pAfCnADydlj4OIK8eipcJ+i6Ecm7ObDUBtF9mFYZM4G3ojU/+h
k1CbW2O4xtUigVfDk6y39dQM0LUDr0zOfOZfuFMuMNP0A+B0VV7x1u0ZodxokM1i
2Pt84EREt5cBCWl3ePhPAdNRhaq82dV3PBbWNlXi4ASMJWZEy+7pqJFrA4deewhp
8FZ2TCC3DN6zdIsJoFOtkHp/O+l3YWFa2nYZ9dM6Uo0eEuWCgEL9uPvhz1q8mgnL
fD6Tros8RJ3+eISKkn1oqqNHUwB+Maoyw+0OHJrl/afbLZN6rfQlBe55vtqm5RhZ
FLmBzEflHgwhzR7iszghqGZ853GmO1jOb/DbrLeRg7R1Ac4wNGRmmMXxNKdUolst
L2Mz8K9fopKAOXNKPfAaK26xm+FcVTul2zxpZgd8A0TOLsLEOUE3xv5NJ+k1HfNy
0Esd9TDUeeuHhzRKZesT1a954/JfLPc8TinBAoVUAZfAnhXGLJWb9HXYGveicMP/
HyPoC8ucS6NqUz4EXAv+Ba0NdnnYjZKIvGrw2Ph+QCx7bVbynRBQu8J001URwYKY
mil/CK9wEV24BdIw5iR3YEXxrBhmK0NIQxRzbn1C65FEcaVYANA2sC2gzQABzvhg
inxFdADi1pCHbPDUEA7RsYXUSYfnbn1LXT6+yTZeff7sOPQ9IiMiQVQT4vr54Mb3
umwxol2TBA7p0F63XGi0n2SU6T+6XGeRXmHN6dGYzTIcThzrLENvaH3hlRY+BrcM
u8S+SVhtqyNnJvGjWQ95d9Ukdv5wfILAsgproLo9oifb30C01a5lwixF/euKFDB6
Gh2s4Lzy40e85zsD8IFlZnq09G8u6TkkI4dg3TvRnbZtECEJDOYVXQJMyD6wH8u/
zHnIUtD8kyYKBtath6NrCihnZ5CqTyVXMlgX38KHx8YCb/7dhl0g37kaDd8ywP1I
LkYPdb8qO5iOo1BvChTSCDqxI9hOXBPAUfPihTlqQDQeedfB4drDMP66f4LkWbZV
xPScut+0m9eUTABoB2tm2NNUFCjrSfyzOIcuNT8MSGQF/B+g0CcvM/KvggbvRM1I
UnnsFaGcZeBQYgK5H45qfY+BAywbHiJi+QZzYkZuyDYtul8+up5CugSbPVSNbgPm
I6Yd8QNX0qW2BwKrr1fAuDKl3SKUBae5OxuOVl4XGmm4B486Y3tcFg7PfsSvNDAh
Uf8iVMIy3JcmY0og72Zy+QvoJoIVYghjqeVqUF75jEM3KMEJ0zYhz5Cl6Xvely6C
6RAim/mzZ/6m4Cfj96dMkpAvjpyOevEa3Nrh0ZdpvDzdKfZLHB25/s2kGA7Lnzvx
yoghBEj+rThpcb6VbL9oh/aAdNdkvZCcizEE0BfF12LwGXmUftg8C3TtlYrCE6GW
ow7UnkJO+BCD5HvGRBvWHMbpUNdHqUPPAOEUEqbhXi/Edwr8tkJ1wH+M6wp+C6fb
/yKcokve4eafwJ7AsIxY+lbNMtINrM5ZEsZ2aqtcXAFc5XLyMGHpOD5hcPfZk+nX
hF/NLE9AxFShlKIni0wBFdkMrvy9UHSQAbhCBQgdvvLGl4i51kBIRLW32g12nUnA
i+TO9rm8rFne4ggT1f2kTphaWZEAH2puiQ+uJ5CRRmlQI2JnVATM/SLo0hUcZlsk
rbEO3HUBk4+U3UX27ktx8c7cSWq2zPXuvL+6eXg8x2jO4FbriydzlI3GNnHfOgir
hseIRoM4niZubKObY5hrOO8Mb5/34YGdaYhPuLzImSGmfFLJD8WJLb4SM9OzNX4s
fcj6Prq+LgZ7B0pnIII5QTyra+LHQEyHdHaKv/Kt9i2BsNVgNwUyQw2XgH+KQ0Yp
M94x314WBuL8JTYktH/jh/6RQT1CZrpq8YRA5DbUHsSS2WSC3mBLfnYyj7qPQkcz
uR8DtOTOt+wfn767H5/AQ9zHy0af7U8JPB6JjR1i0WtYG/nfpWzim+TM80sbuFXH
yOlHFg6Juh78Bvf6j0lJAGooPggXBrTgMp0Gjs5wXH0tG1gazQHPss376u4RJKYH
yqqMZq2T7maSPzqErOVyWGCa/IEwoaNcORpxGo6+STAdbk2bv0M+dyjt/780gTHz
RlyH/y4I00A15OmpsvwUthVwWXqkxBprDjLWo8G+mZg0ERHRLB5TWNSWWfNPgdyA
IBHXcRtDuUdxAvTUEW8jfKz8pVbqONWqazl8gLVw6WdR4DFQ7gVHimHfDvXRdao7
Czul2fuGqtHHVFcUXPBsKTmzy8gmfEcUQeXicEv+7ZRjxqpW7B1zCN5TmDAux57x
T2m+m0zbjMBFDK1MQIFw9gK5VsZmJPHwqNGKhE155Dm8pfhQ8Z8oL/FzNSAu+E4B
FWqYaEljGoWivzhDavJCb6yLiOtnSZ7CDTPL6qR9Y2t12b4gp2QM1Gev+MFzzyEI
lVLvaVf5C4lDW7MfVeVZC/AcwBY1EdDPsFYG8k8R40JpEW4MwMeIRuDdkh9YTobh
mJqWUh/QbZq7npF24imSQS9gWEWxT94Jezjsubtwwld10k1ib8iopcvWRWImLeRG
Ir5BieKUM+SmMpxaCLkyyQeKPMpzbEy+PQ6DsWr1Yh/BOp2/SsQAGuS1PQ65B0K5
NDckKPzTHIWU1EHDhrpGMXGsflgrktvDd4U3c5vwO2Rbwr8fWp+WSkkmumNA+Z33
U3hI4jxD0mNxrvLGTDEJbDyVGpO/FKxaGH4m1kNjBr9T+VXTphRz1sTTRWPiCNlT
T272AvhQldFkzDVVqGCUuNGKsfVZRoBJhvtV7UBgfHJqZBhGTw5e6xwojLQOuKhe
`protect end_protected
