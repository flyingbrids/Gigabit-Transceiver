`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bbLA0lm1EEI+KqI+Ct8RflvaYMInI8BIwRskGrSKdMLz1F1r0ZmMkRJZTOI29Pbb
jrHtWWTG1o9wQMbsM70I/Fk9y+zuGcshluYhpEt9/U+daW0gd5jGBbiMjsfxUVfo
CI1iKOBCHZJgmKzAPaPvmUfODF4wkA+fGT3Vy4f6Pw1Pc2XJKsnjLkZxq8GWc6L1
jVuGOKMTveZlNuCyItmbwxR+2YMzkHzvOi8tgSHI67Nwa2znek0Xp0pc9tGfkolW
R4qyN8ymAYiIX25GgV/uZCvajXh1d9gNnc1IenKDAkLD6LDNsQYhPbJ51yfy7Beg
gUR+49lxE2IWMMRywJsi9g==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
WRAIiZ9+U3895W6+BmlVj1Q4fDG9I4K7PVCbKXVJbXB0t1SCdbBvQ6Zhpjt6Ms99
qZD3cNmVBW2KyFDR0k+M9tded8H2Py+d51NJRMf9MxsZ9+cwDI+AnUMA5NfS/cKT
ZU9Az/Po+kfhF+JsIbnXd8rI12j7L/LE5vtB+88BxoQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12784 )
`protect data_block
DokmeQ1DBCxTUQMZsJDbiCcilnD+xOhNnNP9Ha01XzdU4J7XXeC4FI0bubJAXMgl
1OQ1EpBpmwIJioZD/Y2w2ji+nGNT8MLNMsIRT5HTQDGr1o+bzn0pBSUps/PJBRDA
eKE4Rd6N9cSt6mIESrT3KD2i+xiC5cCUuTXUJv3bNA0jBk4v76hWuOw8wAltncGX
SJUSWf1xC0t6g4ngUPHkdXAJZCnMRbnaGxne8tcV9NnrB1CdfuHyHCatGwMpXIc5
CtspD0sT/T8ZWcO2r/+H4w9bTDAgzoxKDO1qFOTJcEAOPA1VCKMGwuyoCW+I2bpw
4EXIZNqSb2+S6VP8njCbrNOtEZ5jDnvCUuzFoWKEIAJwW56iSjJbcBNCIS8lJAos
ZI2W7Qf/jLrOSLimFIjt8sBHaEK2Cuj3IXe/8pFDFKmfu1cveh4xFqrZz4O3E2Oe
cE3XEvElNkob9K9LL7PENWMgZK+M/IMcMnNNn5K3gdAPeALLcM7IXv4KhUXzJjkh
TVSrTDen1nD+euGYLlNiJF7bs2tiT6BZ1vmKA/XknjSeUvCWs3JY1jNLVl/Vcm9p
XvGKmRhpyzOGut7KTkpivMIfNmcsxwTJMfF1aLOfPn7uSKl3gGYGg3m1X3eeaEQI
ns3rhn0awm5MRBb3qQ3VKWLHgMoZDFSJ+zh+drjsakzmUXfSbKSOdbKUunKCc80g
kiM3otSxC/ITKSwVCbOx3JBpI9XH8tDdgdf9SLTziBg6kkV3ihHT4U3FWxeaITEx
F/mPWnFE3ZrWCrL0y1D+T8mvOD+TuQpzLUyQ4mhcE4pH2+RHY4Tzpwq5Y46nV1bx
pOGe9dz8QDjiKWyFT2T7krgO9ENsIuzBFKmYAeS/k45KAMZpZKkMypNecysiLgdN
HhT4yV6M3V/F9uncl2AfAjd+O0VKnh/RFQec8bacq+zfv20CRlvJ0re+rEho0RQw
kPVlVo2r4ZUBm0n80nu8kaDHos8GSZW7BbZWH1sxSUliVtnfhdOyYoCiCGAQo+V7
rmGW5PO+wxG7y96yuhiNtkFlxibTOw114rMouUtWB+qfMH6KC/nYFukDDu+bd/Bx
oCQ8rwbBrKXJxRmMWkXT2EE7cbtTMnt4UtzHBAtKwHRL0sK6U0KnHe3NeoB1/258
Lq2AVzGrwjtqX70mqo7l+og+P399BrTjIkUrpvVBe7sMFEVQCzWUE1T7yLcxvYgH
Nt6BzXtI8vClN4fBbspSIfYrSUuUhfQ47tcGhIK+nMbITNFuQ2Z1mWLXw7ry+X1f
PPnicHqOJmxjv+jOhYgReI/59pZyUhLuwZvGkXXiGkblr2RvkrcAjpDLKFpQKigX
hyKd6waN73MCQnat1nWOGObZ7mT1smZzlplbaxbFbOLPCH/9P7jjAZ1bj3k0Ve32
k3k6BYNBZVfF8xc1FfFQ/wxrmhFZJDC6XUZtCUkTKWMlV2eBUyqMv0mOeD5JvLkg
g7rWuE2t7kP0wLSknn0ZcCNCenPcdGQNaPUXlJ7XVqzX0iDclegCpE0JMXxNqKP5
KqI7iCjj5Whkt9beLfbFuJtJJXVEco0W+Ei8JeW9sll7j8rnrAZCkg97TojeqCgG
6nc5RxPp5tmGBLZl5XzMS3iYA+RTNfOPg6peW29KeeSvPdo+HTFO+jbXdmTSuRPD
9YjItdIo4UpmpvdLAxmHdH0TcWPxrf3+27yzaBhrUzh4YUGPNVy72QAKrn2nuNpI
cctAfghfgmyYqZVT1/kONE0HO7v8AJ7ctouORDBBE27dDybsZ0LWfCQG+lLobCOo
AykhhP93cwXW3UROcUth8zSTn5y/C+UFWyEtnLsa88E7SiRN4Its7tG1S/op3EvY
TFgzviH9HChypcKUlBU0HsUZn2liPVaMaI7qWEjn8OTC/WTROdVeUiETWtsEAXaY
VPIZd3JPHE8KE04TaAmNrY7lskaT7ilElITVe7Le26xZR/1+K8OeGzcFkNLWpps+
9eJvA1W2CuUoJo/yYYZvH7CLMrfxzhLSYpE+Ta+ZVOhxis1/p//FyUoNEP4JCabS
N2k9HJhYom7JihHkRfyppX1WF45tkATEIbxFzmA7y38spu//hw8T+mVFF7m0Ftad
+X9zXBAx7qaSXtaE/xQ8qw96MP9JlnHpCZmt0GP6thA90puo50E8jLuofawVJrvi
XMYBldbNej9CoDXMwZD/ojYTjaZuHVwHQq0CPm4g6vJvRIBij5FQiUDN6xcJ1AoL
tGHR92DIfnwL8UPs9o6gHtKqBBt1TvnTqw1bYwab6GB7HBQNf1TvOeIo7udusSgx
AZ0LysQZVM1zWcyQSVM5/n53KtBmUGUJwiA2yZQ5E85m2TVm/437qkEIeYcWXwHX
qIFcQDcAqGNXOj3C0XZSlfxkvRiWuIlM0R2f9qUnhYykqKm6jgeSdbV5MhOItgjl
VlRcSu8rStUPiAA4z8x9ztdvcfq5RbC+yG133qg/DGOeGeGGfZ763IgAGbQ4elWv
9ceDxgxn82LEgg6Ct6QrKTwBj9LZEIKMh3adcwcKyv3hFkZpZ2rl874wiiQTs6PW
YY6uBPPUmE2Y09LmWGYuU6B1KZRbfrDFjRNZx17fyWQ7nJdHrAQ5I2g76GTKHnRa
Z1mN0XK7xD3NtLa7Epek8Tmjw7hXi0ne11hv/PU+IvkbtRmf3SOHM0hZNnlcWsbb
vzNcX5tsfxAoxijTY+3GwDeZIpTT3XxB3/90ZhNIi7joSJJrz4QhaYXLcPgAruol
r1wVPfD5Bpg/RMW0ktG7I/l1N04vfx38V3c+gFmexvgo4+52S68CR1F19zrzrOJ7
NnDNKlbffHlDIt05ibnWM91CiwSP7gFMIdxUUmcNJsaw6/43nMsU2uhcN5QOdeLR
2QoclbDCP/eUu1axCOaSUT6mfLpan3KovZ4cswKvq+cEU6GZEapOUCnslpHDYlHY
E9mYmc2mrNLcugJBQbswxOAs+mEC0pzHB4PoWroWNLM8zb25Uqhi1LoX1hltC5UH
IAwt0HqLh4PjIGifAE3Xw0f7VtBMqiZGAkUuXmFlChA77KRLRZREvJhD/dXI1Ig1
4dX4S5VdpJDay23PUyQKe9izkdo2FLHuhUuHDL9VXgOGlXLvqMcYSbFX2rj98FDs
lPiQrgWclo3OqsvQVFf4z8i5pMjRDpg6TNLThUSXwMtGwAbuzQXoQEdCp+un1Iww
gHQ9liB3Plnr87r85lttk0tN5mkKp/GZyLBt+aSu6+SXSkkj0GW5J4SzJ2TqzsiO
T8qJrAC/diSbWRESX81HrEFHzBIIug02lnDIxPcxAysgXd8Td9Vj9PAmjwhxI8Il
YXzTum/oUXn3HhIeUzfIRNymJHOKamdT2VBDSjXUcvSk2MRB3oZhRb9qywzAyYNF
oHld40WxsrP1vr2iAhP/TsEnByJmbDyzEKNhBuQEIh8w6aEs21PMrUruW/9u4oWH
XZwwlsIal50VSYDIFWwUFigbpDKUa4417Oq34BFP3+F+16PC/LlbKdKitZ8r8QyT
H7ZJccduoeACXFyg5V9bPmpkiak+h+vx5yHTY2roAs6VtOUfNbpXqmHREkZZIon0
IZppGn0aD6/tStPW51PHdKhkhSG1QVFAC0bxXFrLWvQNFtBo/edqigvdSIQ8W9TT
8W++8qmPLE9XHdwTMOO/q/tkpzvNpDiMlJrvNpxZBVrAktzG9Ae7nElzh0CqF1mH
X1087JwLdytddStPYO+4J2tUztFxqXLdA6QspjRWySwMjGose3ArU6n5Nklkifb9
1PyXIrOg5Sw0U5TjREUGGmAhhxwZyDB2A+nUlz4jik1Up5rZRSe+BeNmiZ026LKY
ZXA+o8CeLI+EZEVE/Us2SPhErpKYDFG+0RrOCH1+fMNzi3KwuhPElmpnPcA0tzk9
4+9nYScDwqaIOOsj+CnK6FgJhFUPH6Ko6lXRpXXkUuHv2EpJI93oOWU0eGI5jFdi
KLpEpId7VL1jajmYPvsZMW2hYmU3+rNmq5FtkGDyHMC4DFiaBvton8JXz/XdqLBD
sHD1sQKutetl5VV8yOd4nsgrJa1aKtcJt5LTy4Lc/npqbTCyKbn8hUltaUdllfU9
p8mpEUzKurBoV/NTah49z3ALsNvaA2M0NqBjq9g/LCxyaUUJ1Cra6J4jT9+XnyqJ
o3JVBd62Q7tiYtVZtzVnvuSey2aeN+VYrxKvUtFq4PU3iDDlB8YwSyhDkTxJuUvk
XjmosXm7C5fk7M17PB1SAXL5ALJN0RAoKIPHBYfGNOHEQG6OqbSQZWh1oFuc9Td8
vB6Xb7E9yyZtTqVaZG1Pja53PZBNiYNPWddNSSZkMXfWsoYdHuq2LnpKFDU3gYU1
r/xoCG7z6QMrbHxXQtn5o0HmKVZX7uQxrHBgJOqyxZhx9Z+MaD6Y/stlykLtUTnY
khTSmcYjNFac/0YmmMVxrjt9uZxX8wS/boayTsZ6yHhXVlHJzh60usESnUQLzgOD
M6C1vg7GQjJoi62qCM+D2054dOhxzZj/VVQ3LsBCNUttq8rtpgGo2cyb7tuwZUyl
hWrsHENzv5VU7Jwc/r582z5LKKox0V42ZBAhRPZZW8uds5EwTHfVCt2NH30Ox5dD
fpWRaAbAVAPiHQlFgJeXUq+LS3FmmJgYP9gM23Jx/XhEiG1HuWsIrgFGHSKo4W8R
Izd6SZ6F16HU0IdGj26M56KOuvX0SCF5Opwtz4X+XTUxAxqM7K6fgQef1HxQbkl0
vXn01sv5fvrW/0TyjLj+YkFq+yrxbU3BD5VrxCSmYFZJ2+/x4Upj7EYUqgFCFMaJ
+NLAulVcT8g/QRBd/h/NzLSeqoP9ewc7/JZPMuHioRhWXpH6E1bFsalW+M93ZXR8
c7p536XFbfZEQ1wBXUWV0IcccCVF63+ytQaPeqvP3B287JunFi47++HgNNKYRe7H
YXqUgaP8otnytlMOQHYSGufUmrb6aelG9jJzWaSAfhdPybevsmAMuRUYVZvqhrB+
O/w8qWTm5yrPlBVU88hhgz9z1EfF2PhTN7ScC3BElbKqaNykjvpkuNSX6HCFCc8c
/5l1zCk0aiOovsMVi9vYJvRhBoQwzAQYRRf2W9ck2k/SUCcPXmElB+b1ODZq45ra
XpBs24FRnm7Vl6vdc2irIZkwE55a98NGaq+umw0vpjjENob/v8oNQP2EMjCtPo3T
fYw3gA0IkrsVYsx4tyXgbVuYu8kFitmXbtkMuVw46Tms5i/FU4WLzxcsX7C63C0z
7m7UTGcGpHHQd0kvTlwoqGk4k+sg+llH8CSDYG+QeGhTeVHPVPAYzDjDW2hUwHV6
h3dRR2vzgDA9Cx4r37pdUS3uDCtSc5BO/1PHaL+mIHB4Xa0HOmM7mEBXlZEovWil
k70e0WBR2BllxgzD7yORMGe8OBsyEtgVmDP2fJGcu4qJILHwHbPvFsnubMaTvnrC
ezSWPFo7jVg4B8NNaMTqlSwtmTGPU+mDeh8TIInS697u2Q71o0W95XSU0gYn5w/d
JLvwyvMAA3e4a0Lw5AclJubWyP8kcydWtyriPcaxD1Gy0qosVHTTQXTp06ucy4qw
z5oLVPh4JO3sPY2OVHhN1QC4Z5qyMsNlUx3k0Il1maJfF9chQklxUvONEu48g9V1
UjI6KoeuGys7RI8j6/Q5IjM+qvRJRQf8eZXPL2q14+KXp59Pv5x3X95rTG4SifVu
PhLjsV/Lj5eYNCSYk4Yje5zePZsr+rpNvRwnioJrKUxqzu7A0zOpmSHmW1q+U9q0
klSB17Yquo1dP4L8ccyqxybN0rNTvBX6/Np7R1wtULRjYD4QuJ1sdaM2Df9y8peB
vOa8EZ7H+E73eAYd0SQFMgjOxgbC84Pn2/mDz1qfM4EdVdLYTmAZzXQ7eDTiX/5M
e18Z9UzKJ6P5zi2FcHOsg6RrPJTNPY8EhAd6zAUKwTjtM9x/6btFanEUGs7D4MQn
8vqh6ScSJV2+gMpb1KMcUH9TyCuEMOi2I28IP8fiq3V93vpylAFMFVLNGgNCjDfQ
jJHuEZ2T1Xpx/JMkbH12kBY3q5gUaPj2ZZAvQQBPErbK22KFCCbRfRyZxIUge0TK
n3s2Rri3wT6mWP2R4bZ9rz38OjrDcmAcZK1yiFOJIXVjdWULoCQa3GYNMRTr5ZPj
FOGlTJFTtk1ntqMd5KWYFjWXVoQ8l9MRoe3OqTfLDYA7L+rXIdM4EESNs7+SwAEj
wxKn+ssiDi1gRnHuqfh4k9kfWYbQyiBG6NKrcUlgxg9ujd2NstVa5PVe1X89NUG0
tFVuj6Z5JmJui06Jy8yEEqj1odhQBjsRIu4C8vJRX01L6dWy8OzdTo8UBplr/Twz
A+71fNGNcOm2M1YC5aNgyYYlI9PnfJQmSbBqx5M6r4IxgGpK3XQS98awhqCXgbAy
aMRxsCH3DzXLXII4LWkdB2Qz05G5Ds2zaSNWfh3/RMKmAhxZ41fphgYKULgPgqFs
9cdZjYpKtxO/VS8YeL35ZpQNaJ0lPN0PDELZN/sdBul3hUfczSCEf0CejzN5D50t
A9XajAGPIo7lqRK+PfygsmRXiCemPEywg+dW8AjbEdjpcagIh+RgSbhP3MILgEu+
d5nv+p7UebY8Ib2Fayzuh7lkgNaO3ePeSunzN67yjUL9am2McGmceM0fszAaoOdq
MSw/tcRnKMVeDFst6My7D5/DPgfLzQzFQ2vTnWRs892A+TTxe5wamU8Ul70QETCj
ZVTHwBlAhhnacPSAStbw71wbD5vIQYRa9Z1Uvzt5AMjAYQLA2jlU+fJzmKOaZe0G
rn5zD2HIXtfJ7guBgyfOwQZ2Rm7j7JVYXSFl4QNmJINJgKOpRE7Y9rOmLvPuGf9Q
+dyJ2QTtcKhU+eCbqV8D9FmSAiKWtlNokfuZTBlU4lLhyyBz5QE9USnJD8ZBsous
GXiSNVKchC7rWg7URqx/bm5GBt95ZaoD7ZEgjeDCaCACMwm42lNhcqiIa+mhaKtK
erCSJFe8oK5U+lEnhcH0vuULEc4fNKV1laD5cKV16UuZW1/h+8cXPiA3IhsJXORV
dPJMmj5Q+5MyPPZ1EjtMSCbJ1wWGI1L2YpDZY8dUkZqD0O9su73/7FtXuveFQrnk
G2f3hVGn4oAa3ouFDhD4hnosKJMrKwQKUbqei+sl02qBwkC2oauwUrSM1eSD5Amo
0ZeCYbun7SYtFxjJNGJbsP/BCvM1Sppb9wJxwNlLpto9TY71P8GUK5tHX/WO/F03
x+WcG+Vx7iWqWfPEbdnIqtVh2GP4bx5eoWQUEhvMMRPoFxFtH7AguFPL+JP4XJSc
YYOD3IR5CdGzFtw9MQQU8z6kfLww6rIiwA+f0ensYhZlESoGHwZ3r1Q9T9ePt7dz
aoJyqNuj8o5vURMRK/TTP7/PHp9RdRxL4jyY8cgKM49vjpLVKfCPHVL2uuNn4RDK
AYTddwoQdRg4RmXHX+VOqFV65JvzL7joRxARngj1FMWFfWBfyrucZrNvF2TMXe47
8XAITNzE6Umuq+8XaQONiSw7wvUg14K2IdVaB/eFqvBMF4yEMsUAHVvlyrccbbq+
RtG+B0MDoaQ8x/7WykDwYeU9wW3GGpTXQKaQlGHq38MC6UpB2rrpfdKU3bYK/Qqx
uJNN8pPH62mpFoso45Z+1p1XEGPnzdj5jxmZ+8zvARnD1LbPla2vkKFNZoZB02uh
So/9CvI0fq9iaegd+5yqco6FwONo31SyG+YN2ncdW8XPJjVrcG4Idu6I8Z7Zhu/n
qcgKEficJpqmZYocL9PtNLBtW/PI0eZ90nB5zWzsz8O9XhOoJx1d003lq/qev3QX
qpISFpGy9zYh+2ilGLLIhZDtnhuiN/Vfx3KDUiviFXaFzRjgQV4heLJ+C5k0PL0p
P2LKmsqHcjs8g7yjjUN8dJxuhoQQKP7T/3F+M5ibzxmlV5YR1rgEqqTFaoLc+dk2
GVeNAe/H6jn6W/dQufEArscRVAnIE5AyefjMI9njW+p2P2v79VxTCh1bQWU2w1dD
7pTdrG3Ud1eOh4SW3eKYO6HZPa2C3kVsCjjmrb6BT+xWPhwuvH6IaHfGq5pttykj
DmylKqogSfX2uXRyyEBFlyRM3fi4J3Q8D5DTK/IJlh4ssl31zhhmbyQpU15qglgT
lkTkNaxMYoC8fL1Pt3pffgZuKdv5tHtTQ0jAXmOIY/qAZD2h5BgmS0p01sAbob+M
6O8cA4l5lWpbHFsvFR/KrYZTvdKZcom6+fGBp94Qd+VBGg69s/kYSlfjaYcCyYCz
GQQTmWKACyEYgQbFXEaseJuccW4su/z72wwK9wywpHRkzfIgTjRmU8yFZstsA4pI
ysCfwUwz07jHufp0dqMyrlDwLEMcDAC/maXvyYohDcaa9jBlAbDjnqUICd3nI1bc
LgXs1sdFUm2kxUN3+ewoK8K8JF3vPXho1UFAa4522Qkshx7FW8ns8ywyPMq8KkIf
rCBrM3hniUiHiTM2evW5ePeHlU3XcqHWnOfmmqIivHIFe/+Kj5/c2UMJL+39Ebtz
rz0nlNX5tiqstEhFTk+xbOFr9flbnRRzKzQZ96upAlpGnAjgF3JIct+vEnMYeiCJ
IPov2v7QhJpbtokpnSsgLohUmKPQYbDjVWkIwNqmrPo3kHEwE6k6mc7ZyUhASNF0
2sQULnzkWGZEymNcZl0mFcoTn9kL4m91i5rNsSzSjMq0MiuGmm6d1REk4lOzpAZj
Isw3qklVAiSQFRlwCnouqghVz+Wbe3meQ9W151ohlGbpQVBTKB22h5tBdkA10fN6
8HuHiX84BOjmyxq2IqU3Yz50se6ovUcUkgotHINAUy3cppsxIylldGE7AX2IYziJ
sG5MwIs54Bh4Aibk9cJ1ZYohlClQM9dOy2DT1o5fDxVAxO1MiDx3V9sbmtsxWkYI
dOc0H3P9nJcBYS7ZQtRso5IM/juufRNhF2x9EFAgdReSpJlV/KxSeTQxJqh+aHg5
AEzkjarxEqb2L1ME0yAO8q6Pdd80Ban3XHtfLmX6MXy7cKINknXxdyZ0jzI6pUGq
4RtfXdQYLwvW2Ic+CL2D9afjnaufxB4EiZe8vNZ3qhiDHuNEQaoN818iJEg0f8J+
q76RGUEOslOqC1WAZ1SN9+fYfPsY3tBIhx5xLKSW+FxBBMgZaIKTQO7oQDxiiJy9
HsyveH4WXmr6qsgyzUelW3s5pYB2E94kDzLCS6YFW80dlpPzqNq1G+kcKR2OWbxo
ooHIsyD1bbL6gmbigGcgqpLZepyuGh6z99wgOR1dTIozirCR9P97KPrhalJ6MqXB
eBXdl002zB/dKPPVInlX6mzL5aFWGVo/+FfdEbiXZpMRp7AhEMKcqVQo7xQVqOSs
xYMRVbEfRtB2we84nqZdwWZnqS6QddpgYtzykpsFH8kH9Bivj9O7mwk6M0TXS7vu
uauQvldWgAoXmvl+h+RL400S86NQ6nmtUtanlmOEOYVJ93vaJXb3paLR2hVcLni5
2fTS/ammrO8SX8L4KgVXDxCnyHBnw84zXVffIiCeINttLvmpApYmIcpSJDnUdjqT
hGB0/THhNwpcg62OB8Khkr6myysen0Yaso4ST0+fYjlIxErqTiX1TpnFKpbI+HlN
uWUIKK47bxX+0T72vxmMDkdgC3O36TR6HrBFmYLFGnfRfQ5nbPZ0+mx5PFgm5CVz
92Ahm7fhWvbgmd29oYMv5rVlFB0/NltB7/SQM9TiWNHRwGsQJ8cMni6yqaz/SPFQ
PKb2UcjXfy8Vbnz25LWoUsCETT9vMuTTO3U2WIMF4z1cP36YFOJ+I5csTxJzLmXi
j4dWpz9vWszJyRt9oNPolkqBxxTDBQCEOmO99nQqdDp5nplt57HG5fxZBbg19Fcq
RUoG+kcZ+Hura8BOFG20tRZPKSLavu72Z9fOvn1tmTUsifYEFkkNr/HZZgohOL4z
lOCbb4mIpeMffPDNr7W3PwDPzNpY2LxK3wHuFF/SHt+S9gasdMHuAPhkXRQ1c1km
lQbHJRPIeDNMv42/lQss47/7hMBpsKTJrzlT4LCgt7dLwL2h33YtcUsnGbl+zmoK
leWDjO4YLHmTwVWp8LsE6znSux7FjXrisKIo6yMRV/tv61iIgWIHdHVYHFbki0b/
puhZe0hytAD/aqVBOwqkNypLV88LIt8jGGoTMVg8Dp3bu0XXr0DXd5WOsG6Q9kqh
IvfDh4C5CHoZh+Z/mma3ufnYouJEV3GCwsweiDCrjpbrbkxFiNmOA0t9qPlLbBJR
eEkDTgG3GtW/qCnN6JlftY64I73MXS4gPhkc4m/K9++x5hsCQZgspi7SARnpunj9
EtgvzVJBOGJVXxisinJ+tws1gfOFD+D+qIG2W40vyQtYZoYWO+TIPKgAEZGTxerO
nJnvbYdKq5wkQSEZTis46DUmFesdr+fHqH7XoSskPX1cGSKDC7QXJr+qV3Fsc2lT
MPTBwnKXGBcb0nXtIc21XzHdrL/eerpA/+W0esYnvmmYp+w9WgXT7AV5wTPPVuwI
mE+zTNkQt960TvmRU1o/+9V9lkWP0+qcTyxMfafpvj4hmvnthRxlm15quVldJqAo
fV4S2Mmmd9SoOtRnJhZktvYHJ4wHUZ2haeU4wNITyjIBzVpfIbNvzvlpmJO8rpzH
8uGn1n9J9cbTJpM2ZrocSIBlddy3cck7qlZVqOdotxFu+0v5Q1oHs/dh9emXZBeh
RrE1JmihISRxv+hc8R3pHW/3h35rdme7jVGqsaDuD1Csi6vLWHXkjMrGUjrKZaNC
+Losv496cKOvalL5hYj3wTRoVLmyq0WwX3ZThLSOG3VELthGMrr8VOJN+CXCqGY3
nijXastiy+rtemHAQL3cz8H9cHZSubZ0CzZOK2rxgUCnC4P5S6xA2fkQcceWPfI6
+VPSdtdSURgBrl/SiwQnYeWTHLSTm8ZbQ2n2hvvHvTtH2IkHrY84Fqfnpi+hABEr
6wBKlKYZvFbqZFs3CTFuZZMUrmzW+qStmscXPCSj53izttubQ3Cfe0KqAJYbzbho
jVxzspKeTo4FohHRdT/yKI5nAMx+ZlQq9Qu2ougnAeYMg2xPbncuTPS4lG1aCR25
+vsEqSKb0c+1ipyNdfdYKdi5VGYPsRIsuoq4OiRqSCCjyUOhmA5YzU/ND46wHcyS
so24R5hCSXsTdq/37atJsE6JpOvJnVI3HCIT4d/7T+ADYtAhg1AjkKF3glOA/oM5
WUA0llPIVU/pGczgNCbr/JhZEiebZ36IjC+LDqc7YlBvdL127S9yhn5CIModF4/5
m5n7S/LF3eOcRgnPENhfik21A0Jsm22A7UaHjiA/xYtXj6TK0rufXHiVNS/dZvo+
17SuDf2r8MEGxXwtt/BxuN5KU6ePaa6PbGf/cE8wAWavq6HFWQLBzA6WcIq+Yt2R
ZmaEL1rxft4dhLU5216OUkzvfycNZ991JtuSgKBIXau6Ylhmm8CQ9210XH3DSLgm
YbEO1JLKkl8+5bQ+wu7m04LYAAWPeGgApDyfZ6JRDDfbrNu9fJRPn/audXsuhwIa
0GJ4L0EHuBSGrxJiA5rUj1xkWfP4Fibcg/rFS1TNwXlzxs7JgB3rigPXanvcObt3
uq8KiM/sepeNBZassAGt6vvUaXxsVHb1NigkLiYy5bHvGwrhuRhomgrjTITzsIGf
vYKAxEtcdApCND5B7VsAl4twIknIH4kODgK/2Pc6sF90yuGhNSXxQF/rK8pSeLFJ
FXInEXVS0+MhdE0+XhO13M/POlYzyjHGoG4aMG469P+cunKj8OYq9MIrQ2Yon48g
TokC14I50BrF0A9XVSW478HzUDmiMJFT9rRSVKsE7Iha9kE47u/ijEXvuL6oZbeF
DkaVJJspgCdluOH22/eFRVtVTXdjD8ck/Chovx3YG/km4feHeH3oQ6xDI4lkQyOW
0uR7CMX/r9V1ZnIqqK5Cr/yrQP495sQuAnmcRt+mPrDlrdgd7JQgE8uROEhKX1a9
AGQ/bnm8b88YZqk5Ji5RXC4iIitcnkh/v0gfZh71zuDGVRa5bHKDclmUn0+IAiXe
5U4x+3JDKV03cL9x1BfKzGqaXNGCWxhUwMk0nrKA5qaEu8rbbUld/J968jMmD9od
gdCHuKfgJR/RVideNVPsGSNmJqUfhd8cuUTn3W4aqzYWD/863K9H7K3IPLLXz1Po
kWPYmmfPwR/+A3Sv0NvDQtmQtllWrbM9BVeqGQ3mvDU/owRybXhzC92xONq/LAEW
O8fIX9E7EuprEBhdCsIDEn0DQrHID++YcGdBAIkm2RyCcMup3rgMrPfsbxvy4GAW
fnnnT5V819aE3kd1v0/fpt+rf57JvO9uwlofSNl+hL7MIzCQ93Dh37ujZ805rV4j
cAU3ZXFwl7O+c00xz7Dl0BXm/4rLRIg4QJyWmYfUL9CmcfI/BlsPX7IwzVc3j8ce
Q3d2DfR35mDNEA6MzpFcKRzz2+HnkUFOXqKs+Glhy/AGQ2TjU80vQ7U38rDWWYhV
L70/hn+c4O2bOdSAO9SpaMm9zX5Nbg9jx/dyskpq6pLCV1KCYeaEbwYj3K9+G7PL
sTr3m6auewYJx8gZxBbRpDH/i6LbCuwJteSpqTYqG7JapukDpFsG3fWbmpclGsSq
DB65/dui15VMDr4HyO82rJKD6zAGX/fnWI01H+rOV4izR3YUX7T5WeVIqf7XJ8Sr
n119KqEhJUxBMV+Ke8O+tjj7/+k973wo1Cxfvx+kaacsUU72yR5T6uqGBVIws9Qt
PnbgeVpvaMSQEXSci2qKZuVoOl9MurGBZ4oLufINpooiGLruLReO+QapbWnGgYTe
lMttYQJvaVJF0fF7jPtl2EJ6OxO+RnCQCFXlrowT5/vobdCEj/Abb/ojKxTrknYw
engoYDh9Cj7MbVQmGtETf/WEMOqusUuOdT/f/1z0txeBgVDNz6+jr1qgDQk8r3Mc
1cThYj4ALThjQUa228QY6vrcRf0Co4Cjf4ZsIXkOaAtrAOoqP/CRYfSgb9SImXXZ
EeCqWJIRX0R0KqgJ5qa66Gf2zpXIaYtmKPvNu0FUFy7s9pw4hi39iA98XF/OfEsz
DzOfyREX9vLBcfSXfL9A+0fPI1dw0S78TMKyCe23oFX/dIjP4iNX8F0c+A5q1e1g
mLGrQf6vE0gJJdLJKAeD21qv1WkSHU/WlS1S8XSt8qtYJx/LZXPi8T3UhwsSQ8I5
HUNhX5XAPutHK1sQi1iFu4uTydhtayli0TuEIL2J9kT4m7Z5XDpa9fXP4hycTO5g
ga8mLIlgdNppjm2qhtzhxKTblVqkDuA64NwpivyBTpBEj7lWJ6tBeaLlPsShAg2k
iiSYyHvF1U9uT1u7CJTpU3ZgXQw3GsPjPU2DbokkVyzPuy3VBlZq4UUm2wT/4rVE
w89RQVbIW9wHhJ5Ybx3XZduKLAAXvFylgquuoxrXiFmHpDFK7AKfQ6DK6E/dm4g2
MQ9JEJi+G6LabUUEb7up5KBJx5gnO1VeczeZIQiLXVI6tyW+SaTQP5KWs2SlMfc8
yo3lsJ280Yklo+lq+zAywOoTL7iaBCm44nyRskVcOpRviTc260mg6ff2P8YeG+dc
LbGCG9gTPIfKyCt7wxvrcd1n8gswKY1lrTb0Jnyr1F0x/XT0Ko+Rwg0XfNdnedXt
VsB9119BtsGFSBb7ao5kubsfJheOrVEx8jWkUNhs8WP+b0lStY/Qgk079UoAmMc+
UmMXsDbPUXr/t6ybLH3iLflqxXsTj89OLk1nX6qmBAB8wZFkBHTl6wQXwF4bF8Wv
6/CUpaPgBmIvBXsI2O2+wHoIBaa7+9xkELMXVwS/PXl/kEqSJcoLHgXc5hXC9SkH
A2t8HxS95bSZ6v9xylLvFPn8R1+wBBsJyIxHrAefIyicjx+Ktckr9lMp5qfCgxBp
zQsALIrFU+4+r5j2sCRVQkDZsU9kCjswoasZTfWdCX6QUldkW6KA3NbayvlZRNmy
sSqblxRQZMIm+pzIo9LdKkgHj/suzFjiKF+llsi8SHmx8BMGTPIrh68hqizRtXSq
/S0jLeMi0x+73aOaTAqUbibpw+argqfZeKyhTkF5fc4rtiObDqSvxzK3QOHxn5+f
5qXvh1PaVQApFmCAySCRsrPg1MeNkqrWnY6lgcsdzG2DkCwhJtOuY74YC4KfUh8x
+dlg987HwN9yHflSAgr8AhM4aM9qEWepRWmA7yVKP6nEOrw/XC9ig1AtcAN4cn3S
IdoozC72z3vvdv1nPcY8uThhbhAjf9Kcqh16MLnicPkoX+wkvTcS8zvXjWYXv0SG
59H9e+ai/P+MZuL4zLdqqIgYpU4S1zWBInX1sA7cMKP4JQE78lHcZfIs2SPXeoOS
NA42m7YL2ZJUCyHQbcdSDxaCJjs8OWV9vjtf01aE6+dmcJMdGX8VVRXWLv7EptGJ
jRQFEPktZFXG4398+PfsFpzsmYJ34AjmUH1X6UFBa02/PxPMfUUQAnnTccfd1kKl
bEMcwgucGV/FX7Xjtx4FYFvcSnURXroUSTeSb7lZoNO9LkuINSH2TQQ2AuDjsGwR
ZvZ8vnvdnPt80DbWOC/UNZTB3Tc5K/b0sAbNQUhjNnDVLY1cxLrNl+H4cStl6OGc
09BqBcM2cgNXXs+Bh8PuifBSpzfct54RO9OhdnrWQYMHhlq/bpPBR3oW07cof8VP
iw4vY4g8xYv8yeuak1rZMB43KFKb3T1jzZo0sjc8l+UQYJKJgTvd8V2FwtNNqHOi
V4ZuTbH8vGzIsSxmIoF/shjoeds7ufCK0y+m37x1vxbUFmNctMYaRAOH3j8nGie/
kFCZ+Et6cd7JvFG4elVVZxkFC/mqnljxxqYa6qUxVhDdY6UTBcdPbclN1th3PgQI
185xOD1lQAzH6pXG75pEpz5gIhJdfZwshY4FRl8ZNhlcgreA+BzH8v7m82b5wfjf
dKSyyX6HXgr7P+9Fo1jplMGOBZKQg9bDrdMhdQeUrYG+KlMly+FUNSJRtBF+yFIZ
07R9xD9LriuoQszDLcvp6JXBqCDOROm4WFOe0cUie+XVgton1M4xrRITLdFsHLCE
yoTWUHAdVFw/yMEBfFZO1XoEXfUxdbrnUtAXldTQ1PBsy4gTry/dsZamPyz3LCOx
yL4AtnARE+v0DpFjaKT/wbcd3QCfY7ibbZSStDufB5AYfRGcneKujWIMOz/ZOtu3
9pbnzk8Bx0VyE/bIKv4UnpsLbKJ5f7Zs1unfLn5BUOKm3Zxc0hw3gvaQYObRjxq2
eCVtpNaePTi7NRRvuIXDdzTSGhUfV82Ucit1374JpUnEzmD559JdvlV2Px2m7a0c
jr9gB1xpW3J74aJTbAAxPL1UznqsVzrGNOd7ri+nI7+HA2rmyLxFV7aO+CwWCcn2
dFE2zb8U/6Hgx46bsd9hrL2IQ4OxOpHPUxSdiFMtUx1ZW3k3sv04mFFUelGNs5ql
F8FEsRZ9F+4V1RgCQZovypEOHKUdPh5YTAAQkais3gINyujPvnERA51xeZrfbxkQ
Vi2E/dMAa4UZcJRkfc8yB7/8DzzJK6XpE6uQMjuk2kf5i84z1+vVZeMTkGvQEeWU
riwYF+lnH5unpyi6/URvM9+SWl4DYiQ3CRJpMJQHupUGxxUL58k6CLd4oMf82E8p
gpHADQrKTCM/xmjcDUnI4AtE0oziXI75FDTMuRFCKJNlFKGhqF3PKEL9Kw6TmZx7
HcnYhKtRkI75trEcWdZgXunb1bpaIbeOSEG6V8b7dnrrJj7y9iR04MU5wKLsMIBT
UAGmD9vV6QFCzggdWN5P+0YuaR16ZBCZHcC7wOT1Jr5iVlngOk8pf744GW8XEiDN
DDau/zCjeJLA5uRLT/gbvkHcTPD2px0IlExlnVfmlF919i1LayM3hpbCWI2OdVHT
2RodW6YZlw51bL1orWMezHIO+qIDhh8Nl6NaesA7T/iu+TwqCYYjJEcKXzLIO1Cp
Wk+gmBkaxR+SyGNiS/R9Tsbsp+utlVLQ4WHaOEujJQpX2ZwPxhZWRH1MwqGX6zfp
qF7qaaYmdzQ1ZTxK/nRceb4U9PQLyR3hLRQMnBqMN2T1GWWrCN7MDjpFxNUQZYx8
iankVNgRSimt5Fj11W6J1zoZCdrdqE43RxcLA1cvBzd7kF9DWsm8E9Ki97+FS3r1
IfA6Ry5Lsh1zEGtrMK5xk8ED/4DrKyHe0HhhxG9P3ZwshWkI+o9zdes9yJtfPYyU
J6bgb5PnoJCbw2k7oG22j4Ibft/HklYBenJK30s3cTHCG+XgKPIJMoUz/IQarovD
gzEGxXN87qwPmYBuKwjzwoenJQ5FoJc/WCy3e+rupLtUvhMv6CygLhIFWtsSDKBu
rExvu8iRM13DsN0h9w7/jhSf7Xv8+dBPrSg73TQImCR7f+XxxrZQUBm8qfrThWxw
lQ0Y8G4us/OInVV+4N960syI9pMcFRf14drECy//XLwTfNN3kBUvNe/5Dqgpr+08
3qHai6AoO21mZD8WbmIx446nGEEvIrtu5N/uKF69Z2aHhaKmsul2Fv3/ytIXMShm
3pHier7M8Jb8puZD6GbrgMKLS70hrWfF/OOp24zC9fu8vhPzJxQthKaa6ktQqTY9
mLCEFkleOR8VoKXihaFDODtIRHf08UXouiDdX7X06tSFO8+Q3R7Vyp2YIXY1OPJl
0Yrn/4JGLOqWoV4G6E11ovWgHH806AAwcGsoc0iGuA7LZW+pRpLaXy+NExQ7a5S6
jFactw15kA7xflviBswmCorDUACZljpiIT3eCcaJcX1seZySkCCT0TcraIfT/T5t
43CEwudnUA5xSQleys2JTUv7E17Pu8NoePFFeNumasLTVQTr+XAMECIvHLZ0rPjR
gl8f4MUOqAWfHq7HZjdupDAAeTh8+Fe4/MCfBYA2pFW0m8l6aO3LNK1hNvB247DM
clz6dSg+Xpx4RCbCAqTIIo/c0wDsGLVuONwi35Z+q1ZoZykULFVMeVRkMGg/2AO2
uA0jj/JkibtlBRssh/83/Z0wG0oFcIe/CXerIdfQs8QUB4PtnLIS+okVrCQ57Smk
GAc7++r/Et11g1+JzHeJaQ==
`protect end_protected
