`protect begin_protected
`protect version = 1
`protect encrypt_agent = "ModelSim" , encrypt_agent_info = "2019.4"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2016_05"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
uzq8xA9w6xkk1BYx9xHk5bBohFggwzcoP/3Nff0JkENniwgRGxPvf4Bm0GxXexOh
ZqayZV86shvYjnPv8oDZPuxjz902hscVJJDry1PyM+PerQ4IEWHuZsTl3M+11hVF
YoXtFQ5YvIyuYm1owvC2leB/mbqQNmK7sOy0EAr6FI2rMo5ePwfP7m8odUWZfbyY
4GD+At9HAz7lw9xucqnNdVGtph1MjHHXyGiMHICjQ3P5arfe8j5aNaBZWE7o30eS
j353Yio1iEh2OXc74G2iqWa7jcuUC3BItQf590W4R8T1GUaIEfO3OG9p12D0Ri8l
FdCvgZS2JxUat4wxurvYfg==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-3"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ml+KkzuSBWNewLsGzi4zw8mS3eYPDGI9GK+njErwNRrPVa0q2CoUer106khaUYnt
Q0q7NAgfZTzV6a3ehXw3/078JBaOQX3x33A/4hZB2obvxMMMw3yiE/q2urfxWC81
Q1cMfEINaEdc6Krb5jhs2+IrE4begKNbW1AQT3yLGJQ=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20112 )
`protect data_block
4IuHoNEns9M8w2HMLDbKoCD0aPB/M92LTQogrynXqmcpL1WnsXOWb00SMpHXw8Hj
DZibyQ98xdesz7KUiyIaHv85uLJsS/ZV3gmrgxm0a5CSnkBWhlVGvgwWeKYJR1Fq
MLj3PQ1wLWq3LeQqH2x4SEf9wTFgyb3Vbx66KUzjHkxiREjcazHQ6vg5jAlhd6w0
CIg9zrzvWu8Ren0pCRPDES7JrU47S6Kr8vSXWvomM6p+4V/koeaGIjqwKinWSjkF
Ien2ZA35Mme3A2niTDjEQphNZ/anRXsh0yTctacg2+xzqjJgrFlMRtnUUz8l8xZj
VWFYKWa3ax7dx1rGKo0G9JnMNuhei7/NNv4S+Xk+Nysg5FnQfaEwEVZ75opY+QG7
Sot095MhvbgaZ+tg8CpAVoq1yOvp/oz3iAHNaXoN3i9t2RfuaBHGmMhZkN3Bs/qH
ATN/gqzeXRmOBo/+cbz06peYZKmPbxG4Y2N8jeJuLdomMRyBqDJGRoRJNbyFUfzT
u7K9VoILTCjx/b1j5vlBlPLAG+Gt3bctaDrw0QWdO6yvPKmPKDr48nKXQUWvJ5BF
tJPX8ARorDgnUXqBFYLJcqXmbcLyIfb2MMB0Pzz6+N6DA2PYPGqAk6oXVMnWB4Lj
MSlsDPZOLtcDIO/zJ4N59rtzlrds2jNoVanPqVRWcVvYJ9h+IdfrHgYUNbT3EWaq
XzN+SRvw3qIEFaP8pnY8wsVrnoH21E0zbIrJ5J7b0HFdLMFSGZ6tEIo/hj/6vlsY
Hq7HFcohTqNGB4qE86J3XAxPQUPImanazKQVuCZejP6w+8722cFJjAb5Sfx5znbo
IEY9ZeNgA258CmIlouaTe38glf6QzzSrrQB4iRkL6LMY0xaww5x6c9J0wbiueaEg
V3WA2exFtX7Eg6+ieq0Uta4WcmMxVbvIimDTEak/YYLrlMnybJrfn5leuHYnbQCj
N71GeU43lE40UNomNRuOhTdDLjFmlTLqFwxLmGdg4sKniSTiRZ81tjYhV9s7HrE+
qtf8N0FbOPqwjCIGx0tgpgduCofVk4nZ/ChajWiplDX5YuiABghoJH+fuOx/MXlW
rnjO1GOfh8J+r41VOu+CHV9XMyaFAxi5I2aUT/JRRGjlynoqzI9f1uy98avpqDuZ
CxGyst7R6uKiwqbjnPWr1PZdankGVfuMppAX0TWCgBz9gtLuAc3gGWEvzghNtOLO
48GVVuokB3WPhthl8uPXpeY/y0oiFUYxQuQ8g51YcKl1gr5xCO/xxl4ZlZLPtzDm
f0gGU25EyUfqXqMtW69hZX/iXhgxoE72U2grszyUgHBTqiCgqZs7p9DKzWNt1lGA
c6cKCR1hCpUnYLDPkrY8gFmQNHoEg/sT9ifep3XCD4uum2AWNY93SJg8ggJ4ibks
z+1n5YaANIwPRkAg7XM0Q5FUHuBZijDE74F5xCmukPu5B5oGJ+cgFqjuvvaOEsIx
+ZEkdYl+f4vNgkrNIL1h8ukDcC1JTTA+e2tZdaPl+yf27GmafuUxVY199IsfIoPF
4dH7KPzFnpttxn/Ne5JwNBvrQd+m8W06JdyLObEi0hMY51LJ+U76stTOvThUbMRG
m9r98bGs+qibFLLrbHutLrsEdyW2h0EKjZu65Fx5vmreEWa+I4+bZeub9LBoJxUm
u6ZIwCLtdFH6kqXeGVA4KHw4F6caB3tLDjnAhybv+n+PfMycLVnrCXZJS1YT1cpa
TaQgoIwVLXDBu8NpRrMz3bNiHzjPrFsv+SOHoD3+GdozOhUw1WsL2iHdc8Ti+mVV
ZBlU/P2VGNpJO4r8qgNmt46lNTT1x4VMR4tP2Xxr1Zrl8oMEPTmNvFyoXPEAnOVL
9nu7oAmbrIJWnBSi4KBqoAKQ6Ooo80o//stcv4r8jlArQw8WwXeyhDfEk+bN4iOO
P75zBUPioybaZM0zWIM6jeapwZMRZEWmpuR+sJqrhelol4Fcnx9rHRi2g7Bz3wr4
sISsjxURJAsdMSuDweRk7wv7OG6nWgRtF8e/PHrM7dliYhWYMueRoIQbZofW58Vx
g4mJ++VABbVHMdFEJYde3gOjHU0PelSDJGSJy53uwpPIyTeXVnXgWz/IFSsA1Wcd
0j7KfObJ1fyjzVNA8q4R7lQZhq9fNuKJx38N8UmJ/sjJPj8HXq68kuFUxCYlDrZE
+8Zw+yusvwAm01oBKm5A/pwjLpqtA/aaunu7Ywa1UH81pI7aL9HJbD7A0TE6E0Ku
9FjG16FtjgTnQ/tiHFqEhtihbRArpBQ0tGQwgmqPdBukNKDpLyId6bzi2GCBFrI8
B/tnyF2uLwhG7CoxvpGdy3xYHnF2ImFUD9xa4HqFDdOe6XfgHdPnKS9M+iifsGUw
U6eQmrEfwUb9gv8mSySUhowi6gSafdQInB0+6BObcfmbuzO5T63GE2lv6L3pmdeZ
XdifoL8olWe95Z0jFFQ0414t5fCgXgMQ89Rk262q3Cb3AiZyYGpgyGi9s5tmrq+3
VJvLjiow5CL+dT7P7To6KMS9nf4nrIZrjf3cTGhZPmTm/jIirposg5O0oIsLc9jk
CSNLd5YA0HK3aIn7xveC+i64nWX92Ka+cK0DxdC3yXc7cb2RKoFIvDam7UdNYwY8
2aPXlyayAF+/kxRB2qEf/BeYUDQWW07GgZn1/tbLXtIxvy6I/fXStvwr1fnEegrW
KhMMWHG3bQ/meI6kku61eVB87uDCskTKZf+PS6E7oVQUDR1tfku2cVa6nb/YLHpK
zCQY5XNksvUm7j88wp29YQ7VP7s72FOJ2lelKMMl6rM2TaUTYmqXoWXC5F7SQxGd
ILaNBAagj93UlVU396W8VioI9iJeMXb3oMehfQCcKafA+41vklzDKpEwJ58af+J1
/7YswCrC1dWzYkJpE/9d6ph7CtbciiLGZWMvKDWMvu1Ywt9XnIIyxYweudvxn8Ag
rHCEJRqqvQ94fM1wIuWnbWOzOG/j107a1iTyR4uxCu9qTZN3lpSFP/Fcfg12VQaq
zQtTn8FigipUDaZMj1jj0vx4aYQpuyk1Dk0BgpF/79C+GJtAW00qMqfET04SPoiu
52mPKKAkoiiZKLLb5GSSqegM5iq3t2/GCEcy0E9bfa3DWa/DXAqhAgpoFId5jODO
ckgdMrg2FMwK6W8EjzqY9VxpoJCKEBejLEQrtUqCh+88eHJvJ8l27MqDBdeV6rJc
xz2nTSkZV8s9EhwsPqsNylvu17AwcqFa2R+Oe7R4E96wEJ0L18xqh2B1LYKoENb7
9aFmp3noQne/8s4gCdZqsfoHRcyOnn4dafk8PKhUsw9B+xrps6cyew+WS+y/IhcK
Sh+4AqaCjLkEGw3rrTS5m4iN27lvimXRml+BXKuifguooYmtl13nV7F6O0u2HS/v
TVoLgCDPlCG+E0JrR4x0oOqSjmHSFGrhAqo/7it+hFFEZhso94ucdjp4y8QNAgkP
OTzzfZUaMSSgXXAg7dlZnaaLN4NkB09Hq3uun9EY+UXjT+nxlq4gEC2NAW3plGi1
FrMbxjXWor/mPMa2Ns4N+AocccPA0DMkKGAIsuMHSruqkQpKbdz8EGKJmJqVpUl7
gEU4mcNgSaQZ5hwbkf9aWmE1oCGDo7FtbXSeoctpDGQj95S52628+e9nayLT2sDe
5WCYI4MNaPj1SXo6EzhLDkPxgbxbnI9IWt8BwcVIPeVh/QH0nRdZ5EC//hGNUvgW
3FaeoFyHhi4zzk9DcE9wuOmd4/1ASG67JglHNeBrzUdENIgy5CQaNfPqxpNyism2
m6f95Y+fY7UqPgM4Ev9qliUtrmtvDi90iRSCvm+xjMm5Scg5fTGg457A0y3O89Za
5P3nIgDeVHuLdGRea3RC9nduBcIa9bkwkrOS9b8h+HkR2AHwbTWazNkWoiYuG76U
DeMSML+Ny/gLrFzfEaEden81PEqMS8tEij7oyxbFD1nGgVsewzQuH3TS2KSV2jZg
kM/gz6GP/JnPg6Nv0aOFXESZX8PDv90xwsL+DTC8wH1iUVxuJXuRCgSXgCH+/2Px
1UOwrnrTomdYeV8t4vmg1+SqQx1rwKSmoIzB1fTMErBu9iyj6q3S2zhpicpoQpxJ
pEaEOuzFnj2qXzxr40OarOB/opApTGRDc7zr32j+krsyeu348ysApMPjWFLT304o
HR0V5V/5IcSQ9P4om+uAUYh/PmB7339hTqXM0ZUiLaBL33QAKpWo+Xml8FxFTvoo
0MRdJUR2n9tyGhm4FneGQqKWKl1GS8zmJ2dRziF05apY0/vr0Y4U9Il6b05ciqTU
WV8XsGMPAKY8d6OjpUWsmiZv8Mn1Ymx2ZOiL+f3Ys9wLCzsTF3F0T5cAg+MoiX5H
rC1KS+UEKYc+aK92TcB/9ESPF04sPV+sbmdvB2N3M+Wj2GDXi+LA5ZCMC15Em4cm
jYNf783MvnnFa7EAy90soWnULlkl7KVSokiDLr3EY0quW6n9e+5W8B6Qoom45bdp
dgp8niiiHqBudTTCTb7tBslIJ7StcqhUR4JPdNDhCpjulFoayVDFD/3r+aU4l1Nm
adB6ecx0QbQCPPdr5dBjofXPK7EMSZlZp2WJFLSkaAKPPirtKf8FN9gKjYaWmSPr
7NAg4HlbUct9xVZleSPIHavwW/aA2SsixbyAQxbL+B+O4AJ+F8FqPBj/5GYqqCmO
rBRyVgEMSK9w0f6RZ9eZaJiiNgC6ew7Kpz0ajpwYslsKXkA531mq+PlKf5ZAzDt8
jUbBw1mWndur8TG3ykT3H1NN9xjhItVM/00bZ7RU8X6En6QdM0MvmfHGAZygAHG0
Y9TtIMKyY+YkK2yVyfVJ1LhLaSXkKaEzeDPj35Xmf/HNnNiovXsraJDU5OQ2hM30
XNPXeuGzek0rNvxYNbYBHagoOayoszesalhiYewrLrvs1nmsIG2eRlUaukqoiv24
n6yUveD1D0IFFRCR92B5ZpzZWNNkveAgNvhxHVjZj1nr3uWSh2g/JnC8BZbQAYTT
tlayzC+K5wKVSIGEZENSoJjhKDKOaTuRjll0A5PXWtZmI2ReFKI/9ixpcj4KRvOh
FGzAzJyWVnP5PsAwiPlYc5i/fVcBUrwFzbcGt8+gT/MZiLp0lR48dY1z5WO6sYSM
Gzr1oyuYS+18YOxJPO59XVJ1rVPZ+SFQrcPrZurHNE+dhtPWzUU7OOZkRm7MjBok
QtYRONcWN+3Y2UYJBEv9pMKrnjo2yuhPqg+tm8OEPC7Jiog4G6TLkrLCF9PFE2MA
WNe3ukssqBiTqnYplg9AEh17aenjOMrFyVxblnt4wezKy6ajTDmBVIStCX5etyEm
rnkEvAUVVEFfII5Ks6RjMRmplrhOBn8ahBCHtVRwsIZnN0DRF9bDJJYt7vRdjgVP
gRDFasoLYI2CrRZiFckpWj/8U/TUdrj7WJxRDxwfTTQsKbEsmZ1EYlTjvNL39yGD
q8QTf0oBH1EnbemAObaUSV7jOhWQnAoggPGLnVHST/5hbiG2q6AEp/0vhGToB28O
xrqeYCDrVE6VwqdLEtMOS1ZYPcF/XLz7SXca0IeQBQnj3UCJDx8smMiLEEp01M1g
az+5mDiu6QcsT2iyY9AE3ckoXMWBAFBR+GNc6hJxOZ8lnFffjoHgy5z3cqlX3VtL
2HEP/bXHFeKha4jaUy8llPm9CiJ0xThKT4mmcaTjimnys4I+F1j2XXbw5hgEKOVr
x7CRcMIzwWTLHQTQwcXlOcKm4W8DZrLVpMMkIiC+bumCnb0FOw/TuzC4Tif+bkoD
u8rIqSoY6pZHYSlow8P5ajkWGo1ckdcKsC4T44sDNkg9jbsYiTuiZ62fIygvGCak
nWkDeas2qKPNqegIM0SJopnk2MHDtG9f9RA+K9NAX91p7UiLV7GTWmLp8GDrvlFY
1XfFYXMi7uGl/fyO6pJAyjhrqZRsnRZACsD7l7f2cCqkoG0lMjNoHux5ftlzK7FN
wto4HDxTXxS6m7Nlbeizy5su+7U0sVGsEkhiwFOmndhYsCNcAlk6cIxlWqelxRwc
FFnGynd6/NKm4HTWwrsrrDfKJeZp0zt3VLlFo2/tAMTq0ECfQbnEIYnF7seCGy3l
9ONNlywsU6tTWZugy1RIoLVELP/4d1vG2sN63zgQZ68FDc2a4L7GKFQAwcuPSNOq
heKWWORbRIfMAjBnT+A83u9HJ863qAFzex7PpCkc+og4ytJzAdgkk9Pk+GA9/5yh
P8JlAXodhhh5wNKQ4KeoLdUHVxUKGMYbeGKROV7PD0mQdmpwXZLCkvPksHXpNZNQ
Ut/Ka9Ndd5fTBWbCJc79eTpXtZTTLhV1kK79TBlqgvxmNaZ0ss572h5/hGEIxruo
jSSjOOmp2xvc7pcyolMX0NSqMa43sk5gHxEWWWnL8zZOFHJkZd7jxEfjQk6xdBvC
elU12klBrVM5fcAvnppjyG+/ejftb05P2UMK7dfMdMQnR32LNLxyUYns9sLVF9V5
M599Z/7r/cWA4uw8p/Bj6oBVFXNFX5gj4tFaDphOVfWRs+2znOpVI7xYxQmVGdj8
6SZ6mqslqs1dcviu7qWtCBso8fLr5pNKhZXQbnB6Xm4cYgpU590vBLTlWUiREOhP
qKnKHdwhm6B6BAErkSPMzrXAK+55iAd5ni1+LKqXCxn/l26/Fs3LJSidYnz7wHvP
0HIzjjSnCQtNYBbyhNlJMpKGDkqKTM1vfwlawrfaVMMQZsKReUMTDS6ZJE8z0kk8
7yfb0X6P+bbtXmYnk6zQvv5TqxSOHQtnVz/MJbhRg7IIWSM21KffB1iWlNKVP8HE
3xvC7YGjQUUubQUdjEG24Jiip+qlP7oUjmbyKRC1XwxzoIC2/hsUFZY8xlFK0wwE
F0RYNTtJ3QZGDd1V5rrvNWA2NsYwvQleQMypTizn04JZwrmM6yg5xXflUs7cH9yy
jY+xFp9QPvn0WZGeFAU8S4zL72ev6BJ2xNmhW7fW+aU1qZ07S+GlaWZ2OcH7WLAo
DvwArEyMAU+jtUIqiUtB1JtN9t/r43m0C5nweDBptQqzZ35q6MtAh0p+svbp/08i
iUbXdUtT9xIrzyUroAWf+5Lz/Wy6wR9r6K+nXGkkaSiC8MUqI8VBHbtK5Oe5abyO
AGtpLNd+IEvWqpO+5eDGN/zoI7ZqG185NZcxLJy4cn3gfFqeJQggwMatqnNh5rmt
gKUxkYHHJHgS44Kt3bG372HK7jQksqNR6ihgacEKeNVpXnvDTSu2FUdr0sASWSdN
XwOezOHaxqtDpfMFb/l1Vch7wBAnlnj1I5oB27r8cByZ7OMjS4GSmyeqDh0akV4s
xRbsNtyJvr3LH9HgvYraO1wNY9LixhoJSvU/Z/kx2e+6EGMfulpSYDRldy5a4SlZ
so3eDlntVEksNYba1wxKtNr4i/MZZrY/N3+Y3fYLwuU/YlenAOrONX11d1ZLutWM
zhx+GqhGPMLGEMgB2xp/i+F+2UBbXZhvzJWS212nL3H+pyihRbqJ81u3O1YIRDns
8WMbNH7g2t4MpiwmYeM3Nygb2HyvwAHM8me9Dt6v+JMhf9AcK0/z2/g2mKkn94Bm
yPG76HCagPgjpZDWgjILywrXeMCUuPjPmLO4r5zPuFnPDQHiCyzSUA/RZBvK5Zht
1o6YU1HQLAN8U7ROBcsvqTaf9NaBI3Cwyue7U5dmdE0/8PPI9SCV16cNOnNYY/0W
ItyB+6PFuyBUaY/+ufBKhkGgJvPl92BvuH6BXUlA3GiVo/XBk1WtNHcNckOqt681
1wrLceRuYAVTB4tRab+1McxVlLEh2Fp3eVYFSWwqzjlpjO3QUlLOKkLXJbq3KZJl
XOrmFHsGLhME1/8ZW3v0b4ZFihrPXROkHu5JblikdRWoEHEcAKehUr5LYX17OlPO
fHFA9Xpevk+E6K7gtbLdyj3WvAyglv5ex1x32eBqWxNfGfFzK61gqp6r7hrRLv+E
OvUdQSxz39mHb85EM0unDW9KqXSHNpgeqQZlQ1XRtkBPH2LB3pCanWSNZRXCWYd/
UiG9/HhqvFy0uA3aQYpGvPbUJzefi7MgpPmyQLJabFYtVHeKTJ+qgwAOjuRRcN14
AU1K17t2/UCFZxGofCiOTN7LnWiQulAUosijXYEd3aS50yYLsv4a2CRGV2Umg9dE
nP4iyMYEsvsjWHXKwQ2iCRkm+jE3cphaA4Fb5tQKVRFgEK8Edscl1NedX/DyLYNz
nIECKn8C9Xuc8R1G20qdZrD6lopGKD4bTIKHUuQ61iS4ZvTeAoshGtEuMEpYCyjj
qKRgLnElN41KF9/2K02ssGEuh5VZg6oHNLwH2CjaOCHkcbXCpC8ftHM7vWtVxt7F
b6xs8shaIWWXejNUq2BccHIhU7eKcs6Ow4AyW030LcwH6hQU0dntAnHGMOVM+WCK
yNZ5croYCJKOpO0fROmVNrLDy9IIn9xaYfGlx6qlqv+uHd9LJt3GDTdavdhcinv9
PTSu71loJF0v+9NmC/HEciPoXlF19VC3f5GhOnFizbh2I0oZeLmbyAA2JIAiO7tt
VkAgcUkKZMvaPqYAd6Gj4j9HQG/+OhaO1f1+rOmYbpYV5AxqHQqX52y2+7Ep8b40
8e6yp9jdBPs+D6uUCQK/dr0THgiJkBzPNupLdBAeLEFo736H/RVYdypBdFblrdxR
fgpHJAz1afGgWe4TOttfIeOKXccpqPS3z3MSGeiQ8gVncFVgMSiFvuOm2GISrWzo
o+aw5ZtPNu8hk/hi8rbBXUy1nxOjCrSL9jUA5l3dQCoN9tbBFnsHCPSnc6rvJ5RY
WOtVrnl49/N/lNs4n13CR1erseTV3CZGUwEluK62eeI8hA1ha7+FEiGfmwne3Uj1
bzYQyHAu9GwSy5i32GiVJvAmwBvGH3OtuoiMKTwoSq61cRjVk1ZA6wWQ6V5ZtSpo
RjBFTxs3sfdG34OjW3WeTT8SkvgmIG/4HdxlxsZzoOSbndWQDYtQrTVxrtnMPM+1
u0HlW5YdnMyW9Yzg0CeLEP/tCljljEaCAWgQIXX0jv2qbA7lOsMLqk5UHE2hFhpL
k/H/vrJY7SV/56skleHUEpQv3Bz1L7jRAi89kehpj2p5YHU/uEJp0qiLHbiBj48L
n2eti9semGZ2AxVuVp6jnd+t6Vlnd8vuYUkMmcmMdq0W+tGftqKTjz2Jzziv5i88
t0mSxNOUwb7I3wgV1OlyEGwPTMoOKijJ5+luLyzWO+YZ+zPeJC9M6Yq3gHj3UUAT
MnGUkhYw2pqwm8ZDcXkkxiiS/BgV+MZvic8cqCLSW9s9ViUGkLmqpjW6wehubsmL
UjMznAQTbs4mdrSxtgXVuXOfridQ+tYT960AhlptobVtZ/C7IdjWYi2nNBZKIKuH
NqD4pdWtJX/ofeBiEnz6XamPjZRT+z/20i9ABn1w3zanZEsCpZdJpNxeN0gauXe2
hmPDSN5xD+2SzVlTy6e8JnJBpmzHP8acQ2zz5VdiEIyMpig+EWWb+duYbLjtf3bh
80RigzY6maEngb31aRtMjCPUHR1vZvQp94kpYMChISJiMtZxU22kGIDsZcN6gFYj
XsN7HTjCZYeLfvi3CpVyyplakCtn/x8susEpz1RYagaISBKKgwlgb2uun9WQirsF
vO7FOTvFtrIb2yd8p6Gb/hFYFacs8rqQNe0xgrb7G4v3RAjjpgibR0kE9WpAyxwG
bBJJq78EjAYj90RZnAOjhzWyUkpHaLnkm+zsCF3p+UoOPwoEm1x+2pIou9lqlhn+
usqMslyU7bVYwEwF9yZ0EDcPcaxRG4JVVlOzzd3KRsg+T/EurpI3RlWvVSDsDf94
vVjJiHZYcvw3/xfXevt4o9Epnf1lWqPiBI0/sub+TS7lyWhlT6bsQeT/Fgue3zFh
iRlnhd4Namo4Un+bz+3mSMVq0lzUSI2AQYHuXWz5DZAI36WZW178aXQ0q0/J3R9+
jYwcDPr8SrXDlkyAQZEeMcscNIkd20S2PwfyP9gnd9I1nXnLicXalcePooojPNQN
SjmPxFm6glCziWna5hb3/XBOWSStWmVFTVFW4sOqZUEXQqOBiomApJVPls8loinS
g5rJGrE8Ym8SQrLInU6mWQ5zPl6BSwkC7NLriHGltod4zRqgRbzIZjfCmSMyT/Ez
K7bTtFkAChykKfky3mFT+fzzQ5RlSJ82HaDFDsCcY+/Vh7U2i+03p85qit8732Cv
baULXNaBRs/QSvedKK6BKkACs1I/bIUBFEliBe04kZAYt+05JG6hsV0WG/dSAKk5
ioMKKboRGvFLwwI71m574oWD5YyrsWOvlpyUKX/NneK778Zh3M4Fuh7PBW/7hdyj
lHVpJl7HYk4OEh3HuWBz7PuNJonIiQcEtghJBLyYB1b0mTKaibH9ympu7LI7g0aB
TCdEwPl3yr9Zlfz1u4bwjO0XMy6BES0PM5CRwR5uCQOovhgWruhjiB+aZxdGTVOl
307ZZSPbYpvMo9Je/8/lkrfFGqCuqj5SC78PoAEb85mNrvD/2R39LMPUiWoDUMDN
cnoc4a1kBHl8dwUJNcyEfw4cEIIOJMyX9ruJzxVWICVuPJDxS4ISAmnLlj8BW82T
KfU47q/dtlc9Ihtmnb/1Y5OxQ7VlWY2B3DtofZ3Jx+hOuzAorqu6doJxRHbHHfyH
qCkQXqWaY+kBELTId5TsVMcxsurIhaE3Mo4rZ1nssBFyPMc7xFeGqD8chhWnJyFv
FC37aZv82wiNgnS37474/D3p5pjUWPihLv1YD79Idj3/9+hZ1p/g3E2RMId3RJR7
fgK4Rt95aO/JjTeH1Gx0FZA8YN5A0xMZ2HW8eHpLQMEzdqtKF6qLCEdQBSd30NdV
8YndBiIgMF35z32KzuCFNpobbnQou7PJfTIxtWxKctDMaCKTgQwhzQGI/RzyDE1q
3GqQLy/QbpCabDXdi63HV6Siiy+iheIB9HgoAOLms6pns9LOm4vJ+7KiysHt58uR
nzzuaIdxWF95A8hsUQNmDoeT/e8goUJMDBF3/OyjTjDYQ+p8hgv7Mmavxra4Me96
hUCXLNVbBXqXPcoDpt+SQBHLmhpl6qnN2nE9oeWYdYDev4EiUnEJ4o4AYZqjZC7h
MLF3WjCwrFaKxjFMvh00q3fiHldaMKD2ifR9aq3GBRObflDLHwHnFLeiYTCXUkJj
qwvlPbRCjKQMWXhvGs3+qtjJL6kR5wXz1is1vCXdx2+fCzQe7fCzMXd6fo0I1sEa
Rtfu4mKq8lfF0JkHBL/+03KJvlPrnrIBawZ2TvNf4iRETlFDTAVaG2Mnof2+wpsn
XvrxiyWuJ6L6ChYw3WkxxXFmw+zsJ+wKau3qudMIQDxm1cTdPZvCd8zKFuzTojT8
5K64ijHzgKw3XJDIMTuk0DjDXHubYVyR8jAK4rTXpByQcdVMA1LXq2cr3RPvSqZF
DeEEqaoWokW0sq6xRCJ1OgS6uk5yal/pr/NZFRmVSk+H8g6ZS8D6qIj/4DMYmyHv
t84Dzq7yOU4WGU8rUK9xvHRBJGSLlsti8Pwdr0D3Dp2IXVdtDo19wnbgMAbcBMEV
7GxrZNDIp8rZwh18Z79roUB58yepVKoc6UeYVDP43+tV2tZ/5Jn1Xdosap3vbdYt
J91O79I1PXPCqEbj9hQKmx+4Y2bqmMi6hTdzVuMaMpLJtvdghTqgo+m4xR3s1Ub2
uCBl103+ZTk4IQAut2rmjBzVTjuWZNiCXvMleQsp8OSGyIOyPd99DIN+jj2VjZ1L
5b1RxIxMks8RUG7dZqfWjpAXB9xCt2Pv8Y3K85lQdeSYc/cY1RNuveXz8/AF0OzV
andhGuXw/saD8FprXjfbVd+NfnL70ekiW1p8U8xgS6go7Yz80QAEv8jhkz4t4n7h
UjXDQ42kcdG+IVbrcwZJXaLl6OWqfxEsFP8hp7+h1k/UBhleHxpGW66n/N26gnFS
PLzrNBeqfWCrFeBfehoCpY0cX0hM4mTJL5EL9v29aFWUn6+5eq9HUI9TWtOWY/KF
r9yjmx5Dmzp66TjXYhVNQTa2Rs4G08hmhT+odWy5CpQEzKfIOf3feiThvT9g7xdq
znolc2eEMfcjoNii3CY9L09MTck182y7SVE8FBGqcFV0yxbvDGx38xNucOTaKMrT
KUu2pWke0KFNF/1Dgt3xTegMAPYKafDwwAImOpWoEOVkhyR+E1bMRKK03sm7z909
loQ3rRs8vrkzOpAOOWZpuHuuyoyuSAFqEcb1CrCWenT7hBxrjt0I6P6hPSIQfAEe
IeMVvGht9EVDItNBWSz2+1Ajfr4bJ4+N4MKTP9J7NzA2/GRluv4I5xWHLyut4Mq1
FKj+wcym8dGkfBcgW1ghqtFJWHd2dy+aXpT/RmoPh9IvSshka8ejYQXxrGWPeE40
rY1YsZ63XZBYfl5U7Ff+DKcd06TKvl4bPZpG7dK1PWKKMHMAbH2DqexOObosWHZa
aSiSEnVOHnngXUrR1mLMj3ZQhZxP1Qs1YCowOT61suUmEa7nMsRkASRqLgthpybw
qToTwmin5hcVMSiHHlEirSO128qS79os3nVrMloDbs9se8Vw2Tllua/784jHk46j
W/b38QUiLaQf5dmJr2uCcM0ND634BN3+zqXDqJ0pjTNAfswZWIKOwDlpkGAo6xTl
sG2YmrhBxDiXkAUkq6sEu+GGnkz4vMwDPU39OHFbsptu6VyR0WY2O/CfQVz+p6Pv
9PbUe5lXMvEetOcA7ie+I4Zyte1HRqMgF4G4IT9a100rA1kBUUueFpdVtHBl0ZNq
iyHisPyIcl8dyPgAEq5oJtU9o5OrTXLjIu6QoeUxXXoA/1y08qvwiJBinqI9PePt
6FCuviZFgkol8fFNMnoKDBOh5s+T1sfH4qjeP2ImPGyCOPokq0JUu1mekf/WDXFA
v0RJZLRBTk0pu69BLHUkWF0/gp1+w+FqljH/MhLingZH+XN4JlA3KtUYPfhJZhqd
3xqUsz3MjNn94/RzSJajQf2ZfPp4aNng5zPlgdNgBT/VmwpKX6/qQj1P5Sx4XgSq
ic97KsMQuAgABaH1jAOsKPG8bInKRKibnD8KNvEPp8cgRM7z4bEksAjdCE2Mo8OY
pEeV0F51qubxTk5Lfn9/MAx9ITClGQaOHmxgxcw8pFZ+KikjaSo8ZB5W84hmnF2g
8dfQ/9YRFCz994NcGqMNdEP7GM7GISkR+uxxDpMhQzhTKFUcDbvjyYwkLf/N55iK
BxZZdz7mZY1PX3I2vEf8h6vvYYJmCYM9csqobTNYcYxFePIfNm1sZePk+zA4favU
e4vgBUlg6Wybygi27KEawg7DpRa4VbhIY8MtB85QYhe6gEbEm3EHW+qGyKki7GvQ
AWlnEW8lm21xvh82FUj+UIyM0eHVjMEzjmWxARBiPreg+ntyHrPBkZ24YYvMkbhk
chfKhdGlo87ZUZFG9wrd/csXY2SzMZmMWZzRpQPogbmZPI/uXDYhNuyVBrEEejVR
VkdCXoVdI6LFr610kiEzJS3LDKsRIQWn0WUQSJqAoroAWHQO2ETYkRUagXEi6t+1
SvjY2eNiQftjcOGS/U304v0doNt/hJuELwR3zqgk3XPanoL0jZ1BwYbBR+87Gp7T
UbcxyXOl+l+Vy6D5Z1ui5WJ2p26RxFH+B6BfcygUlos7Vu1PaQlf2KEv6QF+GMMt
Uan7ttEfSfQbTnwZtkHV6fUphacpEqcA1YvvPRrnB/dZGshpV0igliq9R7jngkFQ
ae3+0M49V/0LQTYMkO9ceNshJoWDO/ajIP0vIqgcZR4g8ZwMIdMaYelKIZrekj7S
OssIlQ4eBp18GOPqfMBS5fjmiCJivnZbyMlBC1TX08MH8rBfmF+K94i4nyYELsGC
jHqlacUPwQ18EU9GB2jT9H5LmmFXrm5BUYbL9deNGIofvw3Y+7tNddJQE8/P7PNf
WajQzB3ix3ZBMYz3xp9/5FO5j9oRF9IVA1R9+UBn1aNM4+gn5oYmFKVEfn5ItmRw
M9FcK7pd6yt0qNJ36RufchuJAEhhPgZkPNkfIGm+gZozvFzxZxrZggR8NvBEoSgZ
STYkNpeMa5SwSWg7bHggoiSyLfQmkDF/1NTaLB/05Nqwm60HU/ljAFbRWSXlLGWs
rnXxGwdBSL1REHDboEQDRS/FcKdD56RC5JNiLQroQq9p5+B6o4L3JJGKjNPHJS2o
c0TXYHub+pyyV4vv+dh66kpSYegXRf5sil4E7climZUYWg31fKtALVi3naqu/Zhr
8ejhL3PZqpyhkdkQo4aso1tf7zSgyq9J8K/QtdK6jF6IkOAMIYIBaqzd/0rH48Ox
HqCGJw1u+yNvduE4DlpQPaEsPqfAcHLG2w8Af3yqjIcAB8In3ekWy1sYAH7PMO9i
NE2AraSW9rs+D5JCzTjjAeuWq96Vo75SauCUpM8dc58+DmnnP2fZ6F7dGWrQZ/2Z
IapUHTXZr+5dssJWlAAP/esFoobus6aDF/CXp9Bgt1ZUAh+QDxsg+d5kZWbCoPCa
oOO/RL0TqpucnAXn+YHJVpGdiZXnV9us+5dCeNoOZMJNozzoNIGBS8B7UyOoC4hT
KwcTBPZEfo1iTDUY9psZ+VCsNHY2+Ry7L252dir8DaGtSzHLq0lk1D3rw/6shpNo
I7HfB2+fYavVItXyd6yZm4g4afwxVhwXiWJVopr9LVd8GNbogGcOt8NIARiRosuq
MAWEz++sSzfxUZE4XvhB1g6FrrCislz/ZdkNynTfjq7JFxTQwL+6gu1IXv9fHstV
mF3eQkMg1UOMzep3ycntU8CA7XgJu5Hg+dUx2QtJQeGkOeANQ4v5DuHJxRH8p5xQ
rA7h43T46isGm40gJ270oOw8hqcFRpQcf+YGPSDJ6Hxt0B6Pq898qJq89js+y3z7
Ed1YvXwoPr0a3Mp9PyAhFzw1FZaPMUFPasDp+BO07H/4y9f8YTEU/7/KNpL1BfDJ
X9o5xpcnQQFZrbGNIGKq+BTd6cakcLLsDxDeDtMl3Dxj82r8nyrJM8R3vUnAplqC
iuK0vrbcJO/FoGsC/tQRVKD1x6jXzJUHRtGii5f/JHoE9dRq8mZAnhuYzMXsfkvN
kHMGnZbIi3tiyUffYeftl0+Id3G+TgKBw/xJ1/57ysqShZrCb1p43SNnVOeY50Va
HSXkN5fVru2dyD7Jgk4osLOaSh+/RQ3NobCdKWJGtUpDYFgCbI9VcKTcVlROBNg9
6Oz6SwNGtlv1dFbvudp/tUGaSJ055kXa+/Ed6NSm1Muo2G4UMuA/chGk7TWsSFFl
K5t3Ncra9vRfBhrSrfl3p9YfoZybZDnhGNDjq2YUorlDFLXFEec79w3aZdRyNPFD
NiTslnu3Q4BkLd1BLiBHCZbfeVnr+rwj04cFac1+F6BkRrBUhh4M+XJE6UPw5o9R
JOvAv3uxYXvpml8J7QDnFMnfsL7VZgQc5uGCNe0NUfR/niB9sw2a58bWsul9viDR
s4zZa/S+k1/y6MiWyggWi8suKKOT/VPLF9IO1Yjck8eq9zDuKFtDHwihLjGiVvtw
EwmQaQ7QgTsTRX+pmhIWP4BaqDSXq+hqiOvW2LY0vgzJi+WffAMFUMJHH1y/J3VK
qW8tt7yUmija97Nve0HWyAbR6aLCABAAyXU1NKp/WmPBc3dDPnzny1P8nNB6GDl1
d7+Thv9ivdvVmS43hqCyTBGJVGY1f+cqRfrEAJsyn9MLzmxixmMCFIvn1AihiTRF
OtlWwOOsyb9cR3ollZ9Op7tUgZpBmpskugOKJhNAWKsrC87JHUgSdPjAFu8nTPXt
2CM7uEO4ZcGjB7dlv1wx/JVgk32G+Y8JNmpC+c00J9v8nIrNSPM3bnraXag8D30Q
SLaL6Ne20i6DjfWb7YN5G5IkiTolIqcFL0fU/D/fH0hsxnhnQI+eqfU2B7jJiCTQ
Bj31CSrh4wH/is0a/mwwVjmwFy5Y/iMvemr+FAC30B2TWG0MHi4VDjazl1S5hlcQ
XvACixuJHOONDDDfD5H6nZVebRUa7sNbugwl5Mi4Cy8fFJxifSMCaj2ggYmFflkN
yLJNpq3J4m04/P44B5jji/5cpZAyMroCezadryiWD8grb24/QcC2YE3E8G4pzphh
t5BF/UP+XAP7TXRrvxOR0oz8vVOx2T1G+nn2QBumnAmFzRrliHwdrB3C1jze8A5i
WDrxZ4sOW2+rVTCngML1dc6zx1Wne06eN/MGRV3S4mOpwR2CpcTvURYTXYFta6Cz
fTiwgyjp+rlrLNpqaCK50Eby4ykTd6B+M/YOe6pYuZ+INKDlUYmlSI+GNLJojf7P
rtpesi8/O7YMXxuPKZsHe/PtkY24AuY7T3dUCowtckf2rrJjNh3VLNFNl7phZr9f
JeMeN0MCjrBJUlL7JNY7VCdSlzFgCzJVMZNz1rSLSV6m3TO1/gx2R8tSjNaPG2nK
nrMzvh5TLLkiJJ561L136vPgIxpIW3R6jrIRkgNfpQMR01ICdb3wT9YYPQ6BIfGC
i0qIARNianl7F9VKzy6djncTaB9zU/gwWZ2J2MsHuKvdpZMkXK6lNeAXfaxHVl7E
6MQFNKTvUu7m0MQYrz5embH3rvJZZTP6OI+clPFeZ4/ELO4RmMyHbtFxou7lunT0
9QUQ/61/gHJfw5H+D1Rvdj0zUZBFr3KGEgVYF0QXm1djTWQYpvVNkjGXXMyhXGms
RNCj1NTRaS7v/S25rWA7qH2ExTg56h2pEe1gmEUxxYDULsKuJqp8OVJ3Y9oVZcmT
lwJcTJ3eqE2eVcXrUYUHi8lzMTT+siLHbgJxcbIacYMBzawb2WUQgvg34lJncZ8F
oR7PrqU235z3Z4iUITjMZImRYr4g0RUt0ise3KzLqq+imWR8mdRA95X43PR/VfR5
iXLvzLuXwl3c24+/nCT80ETh4gzQe9fzY57/EOjmCjyr8d+8y6mnBm9Dz71GP6Ap
RutNUVf9srvQ+749Sl3clFSGWnFfY9zuS7cN1wnWk03tieVwDhvuuserff+xKZvB
y6ft5hHzk0xY9XtXV6ss10P4vQLXph4IyYi8N/FPuWRxfoLZjFnTKBnzT4Zyp1qn
rTnfR+E7pLpK4Z7DxGJZeOnSHZTv8oQVzAa5XRY9ivVpUr670W4ttnLNpm6yQoZn
FnEESjuJzYPfAnlEnInn0hqSNLQQciBK9lx4tZ7BW9lmPbQIuEqh7Q0Nfevg8a5v
Zz0RaqggqydTr4VncF9NUQWOL6ZndJIjgQY8ZdWUKmoW6b5jto/uEEWUwmrUMSrk
DR40k0gRKKiXbJ0N+xyl9+cgMrVThYAZ4z2abN++INcQZUZcHK20xwXxhCA9V/KX
jx322gJOJr4Q8/TqXbdLIwCd5OdFjXoh84vUkOpR/6bHC4gP40yG+Rr8ev6H86V4
/otnCqhhlJHTflzm+px+ktOJO6WsrHSfakgWGvT2BPd3lsLpsBNeD+2b8oRbp5Jv
wAC2EOVoMpRhSrWnFz6mEYOUVc+s5XtYGL7dksdMJskKrnZA15jaPDQhyJ7nNvjj
vpO0w1KEjKVNq/kYu3lnVaY5hZEDnc1ac0TiJmTCqjrvq+64dMJCpXyrRN2yk8Ji
hNGp6T16RB3E8zPEpCCE8yuEIN1AjPL0H4wt951LRX1Lfj2e9wm3cH88uNEp8Ch5
cg0TUkTEFerYMsFZ/Ieg7IugyWZrO8qGnQNf/CGerLG/Xg5KdHc4pKVy2yZYxcMK
jOQC/E9lJu31pmcpyfatn1cXkVrUdM3lVd8/SBqb/BBSAPmhtCS2SyZABMZddqk0
i/ITS1RuwdNfpNjtGcWiqb0uNcBmHmdNJQwhxTUtdwzKDGNbLQaAA+vegJOLPrVQ
gkbFIBmUrF+aPsyp9ua3pK6AJ0aRGoyq9/Ot9JdJv5XHenh6rZcuGg3dniI2OSrL
Xif/L/49GakHG/K2u9Z9l17t9i2Ab0kqce5rCGI0YbBeCSBHiSoSvDTfK7sWAgl+
4CnCf9OpcOSgqHmJ8UxvstbE9oEIKAAG+BNxqazF8x1MgmgynzFP2R2/kC2R6zJV
QStg819BmNDXw0UJK/GodXVwQ0dXqqItHM4Gk3MyyVjvj2ns8UNnKBAo6niTjY1i
vcYAbeGfx8LE475E4V/KdJAs5lMapcBIIoGhbA8KJWT6tBolOMUe9ge6ZNUXJquf
/cBSmbmgNC/C5fUrUHzjtRQNt7vBiypa3aOeibo3ar9FEF8cyxqkTR9v1x1Ro19D
PwHiFT16avj9xrCv9ogkZW//+Ttg3pbL/k1YQCj717OxLJ17s6euYk1coEj+K+6+
PxznfvvWkFwcZcXVJMBFMOSd7yj20OGHGxw+W/Ukd5Fk6BwbPUvK1oNibYyNe5iq
tt0iAhox9IFSa6SVHKkUNAiUyWLBYgITmr+PMwPqQqiLOGKyQWQi/sXV5azYRWTN
Yygu8apvNlz2UJN1+4lEnBd1KDHLmwqgmuJet3Q6B/ic03FvmqsWA8Z/ozuoOiUw
JDQ8ZV2FC527W15fIZTvTyN1EVH4GDwXGwwPjgOpvhETPHKaWm0tI3ReTNwVD1Uo
c4YkYj+0fqdMDVhVWeGseMBKFrGdvEAYCCauuE2QFPIpSU9PBaKMcpI+qQKuqNK3
TAP+O6oup8tb4qF7UZYlS/l+E3dplgQSS/K7gV/XzL/GQHtFQEiNriUkGud4dAb1
6wPCduibpnbMw7BwJGqWb1AAb36lavfss2MYfwDrBxXmyuoHCyiPki3+G2rvojlZ
rl3aHYo8sChfo0MFmiF/Hbj/uw4T0GNhdZ2t2B8liT4htRRMK19AHv2fXGQmGnGM
UgW9WjRizflf3GmeZ9NKwiio7/kHReHi6gjdMIRcck+6ffhVZ0WjRIl2EeeD8r/V
VwV/l+62XnN2phYj7leQEhe1HVz3PfzamUBunMRbWiA1Zkxoqdoo1qC4KFq0YzN1
Ml/1Fu4EWkqczdmupnhf+OQmsniRi7zanS/caGc7XelGB8CzBO/c77IiWEan3JUE
t62bOi19ocic41/4qpPbZX74TFRZUhomsLEfwljWfVNgQlFHs0KBF0fJD6HtIk/w
q3K8ofMI8gL+ImFJAdkpa3iingZS/m+beh2WQ0lyqbCXtAC0eolJxDZ6bA/mhdmc
kg2IxkWOQPtkuq7zqfobi+78sS44VOM1bDFRTbAOglDpb0GUuQgUK8pxuT3+V3hb
H+6zMQ2ZMBJSDRc6EXowDiWwpYpJ3Jn2l1tbmlI8OwyCzwKziF3a00gQ+3woXa6f
Avb+GOkX3Ih0klO4wMplVmp/fgMGI6xIL0IOZuxZ6XbH6wrYpUTUqtnqhae5W2Fl
QDM61Pq1h8n8tWHFAlC5tHgWwy0Xct6XKgEHeSuAAMcg2PKfqx3qY/dUET6d7fUn
oISTGSt3HRMzCII9qSxU3ZaTJm+ZEL9YHNVNsdaEsXRWjvdPx5wCmEEf82F69JQr
UiicLLiLdUjhIYGii+L5OulFk/wn6/d2AC8VcpzqSDKshso15FTT5nqeAGtCYL8i
h9eHF4tZChnuhN4mtZ1OtSP749jgvFC4XLwox8rH/zLKf4dIruosoTDwHiITmnra
1hrPENDRp+dBqQnF/gicdMXnKaHVogQxChJKE58oXJzHMOm4x2FDJT7+ZeAmyULT
7luPXirtRiu5oFYJ30FJs4NiMQMP27h/ksdqdK6pT1SDyts06LzH3Ni+dZ9nVw2L
yrLj7VFmBg3hGdzJ/HQQEdrBblMdNh//OExV/cHoCO0Mve4vHF6mfP8SLTFr4XeL
gLNu/hkw99dz4K4/Xyh7+InbGUy+E8w+IoXsut5NcC47+/6Ju6A72Ha6QMVZ6EZz
PtvtOIJDDKfNQk1F0ESBggoIJJnfdrhXs0CksczeBNppYOraB+TVtl91dmMMtmHF
ZCCNnksxoicpSnEi8mDdGiQubuIlhZXkS7aIhFwjKlu/RDtMl5Vz0dh3Nb27qazj
LzOsFHCb7Kb/BYC17igFAKDoVv3t1bp5G9YTLh0SHH9/a6XBA+AE6lFJxFq4pe1N
Ov689nNjLM4hpH3DdZk4ZelRkdzPaqM75QVgnDq81pAoe581nrUdrQZ1Mm5/AD3y
0GMDP+hXe9MNzNa5i7BYQVOWtkoudFgtVhTpIjztDrxQC+IwOh2eMV2ZJD6G7/9k
6vW4sPck1XRCwUxC8XypDDtVNK/hM9bhTY14fP7P9COZ5Q/G8U1IK/EivW/VAN8j
4IJG+99xDChVzsxtr1B7OjKNmjhT5hYYLWapWxU13mDy+U0cuphpyR4KpAiO0M30
jlPU1kfgFELRXMg0vaD8s9Jq10HgLjXDwoBGrBJVDdJWw2YieE6jyvYTzDXWEjbX
eC+J7wYTlnM23mjqQ1JlgIiEoRBNm4u3rhUPRnjpF+TjLLSQ4l74I/LBLNjQOIRq
KGbIGkJmWObh/1FIWjsVdIu1CrYh9vwJAna2N6QO7RjoM334STKaKl2XMq+ZrFom
/Uv38+085lK6h5Fx0MTDgFl9gDxuylV1w3z6utv8VQAEpzFtzql2WjcCh+k6DDqF
mm+1GPL1bUs1AsCBNgPgQ7tDZQmibP+FcA9JLLq5rqs9zVTEulByUPBAFIqQY84c
fh/E4pbS8xB1BNxONjlSd9QVdLFBHp1oFY87TndeVdsQWzJ/H0utmfjXVubiobNC
hf75HX6n+RtT/6PFH4Ia/sfAYX9XyAEMH3XRiDOm5Xwsoooje2db+8C3GHTsEUdj
LcmP5GdVnXmNNmVtP9vAzYgKGfk0ddPXyu+StVZUYutyw0YUIhaGl63uuBQTzPPT
XqjevCqqZPpi7dcbhHOa/HwAstwaTROmTzSErnAWZsrVCd7rzzmcxUYk16aOvf4F
aH6f8a4khy7HtiHXrFjfU2y4qVWktFLFYMMogWQp3s/d+qeoD3QUg/5xp6y8dre4
6adEoTvtVqSbl8C5CVqyfhfOu8h/fZNTk+MGYTVtayuNbCKsFL88zmz7FBWuyoQX
HTYsnHxZgs9Qhr0XtfLtWhKeawH6OY6WushUag2gJU585QBqXcY7Kv3CPbnC+ZS0
DedH8XNcGayYAwS4j59H+Jm/os2/3ttSAyKGQgtK00jbbNgHm6hciWxN2jC1Mr+j
wh3PZ3bAbOA9kh9OBjy8+kF8OnNGtxjrRwTMUxSMWfm/VFcjWDvwFwrmnYo7+UTI
ZhTGIcGNHXkSUHRQqo5cSnav+UFCmenYmjV8y14+ld6aTrINNkrGduo959X9FEYD
GjSJyDikxF1oCpYTg2sNPMCMYcyI2l+nQ2QLKRrMEs8IgkZGkzuV/MjH+pNJA0cD
Xbd29jSWszxUDjpIys2iC3EuoqEAcPuf2Q5/eEhquWvPbVCpOcskLE1LL+Q9mBLi
UDYlXWkiee82o7buw6WbjSkrJYTkC/XbeguBNxvsqstWHhQKsYbWEv9C9BPC7K1n
yIBplgwlzH+hGQHVDHe8nbom6C2JeprPVVdzghQ7f0V+rRTCZRTB1DtreThGSYTD
xnTWmbQMNjLE6C5MoN9q7itPjDiYp/HGwJlthGcuWgfWeacwYBeGwPMbb+D/iNL+
Da7pTZtrKddXYNkQAJXJwdvuTigPsBisX7ysV/KP0CVDA3h9YZJppw1ziLIjDhE6
zBxwDkhSO2mLm+h+j2sYTp5C4kE2SOp6mioR6LveEuZyqZF33ZifWjWyx/8TVHZi
+1dzQgcerdNFHMJTStSu0U8xDxXSsDe+/SuN9kY5IvcDt3+4Ipyr60cHF3pRt08r
ClMRbYkAPbmSYZKAINq/sn8WwSRZLI79qL2a8tV5NtuyFORwixHmUq30Qa7NhJfP
2DHkXJnsPGC67XCWpxSNyTfH7uyNckWngO3IRuCJTBl2vpbcDqNFfHxxebahN+md
tKPlG3r1lrXAIiNtRl7q8ihnHZPaXRHon07EnmqrRolbPvBNFQjpCPHV29aRyXUa
OwuDUe/ArGCbG9F9opH3/1zxpAuSjeRThaAFtkSdSB95bKGCpjqSP0sB6i1nskV1
Of5lSvnqkNb2gPO2FC3wLZPxgOrUnoedO8TOGgctCEo8WsbVHn9GHqMDVrwL/CKM
09hXV4q9e1D53qUUBeGS4g9utkRqnwA9C+ncCsLSbrHDY5GsEtQ8UBJpLT+99jIv
IYSYIxGX3QOxF+z923d9xfSj25JmNZvAmP9lxs3E+a2Oym7UzYS6pnM8NuZAoMzo
QOz0tnwvQTp1KxW0d3av+e4qTP4JE+92cpMQ/pKsCAwNNxiTykS/ockjbUqHTFKs
LwmFBmrFmroxnv1jNVTYB/zSNORTGq70N1fXOSUZqMeW4kDkgZDUZAfHEE8nKhj8
WcIGPbSdusUfEJKOZbdrlPYn5BebQSE+1u4Oi3s7lLVqTvw/Inv+MHT7zG042/5N
4NYQRRSLYm3m1p3C0ZaVocxv38CAhKiT0fv+d61kUN9cJYWToeOyw1rlFNaPfYQB
dL3GAt6EQLR4NO2y4Jz4Y3slGdNhaDp6OLGjA7Gm/4ehDrb8knNp48fvjqphAXrW
iLxr67CSucjDDudZLvpY51VGRsyEQbscodW/fOLKz2wKSVvZp3LbOcb86+3SoKpl
I6qhAhAGuzzRTCQZBE7M3CWRSnZcy2+WtnLdEfKhX47rc1rkcSBOD4up3/mOeExL
otEF6by0IM6A4ltg4VD0XPV5Tc06JvXTMjUVpU6mb7u3S6hXeQ9sHyc7ocxdKDvr
q2fGaNAp9JuIhnGBTZ8uj2B99nFHNe9cI9e+RPi3S7X/GmTBwmzbBvaGZqgwVNGB
U4F+cSx5TaQD6nKwPaLt8of3tCNgawHvznHoGIjacmCheIpwTy2uy4lqYbzM4LxP
N6a0ARdtDGc6PByohg82v0HtBrV4BuOxp06YpkcuMmduHoOHkMw6Mw5wIxsj7Hbf
6CzRjQxh85waJvRq77q1tqO8npzo18B5W1Lf5EDvgIHs+BV/+cpJJMuJsVpq1g8b
CtmO1RSVOEOzAyNjWq14HeTEz3WFjZ1s1gEDURsiQXFtl2vUoh8Pgbfif3uSDy5r
8QV+hdWX/9UxXFiObVgRT9zSwvsMYYN162e5OOno6dpVMlhoQ5om1guy5yAuihX0
HZfwRoifbgMrIHq5y/oNIDEvqg5sDb2/vBnGnqmwYd93bUYZG2Xbq/xF+KOLWGFo
VFREWzlxeiXmQIFRhUbjrJwqBYWi3sS3cdPUk/ZezJ9b/s5j3EzvHVpbeW302RS8
5SMBKRhyn+D6g/xaK5foteawAO7HJ1dwTOhYsACvCTm3IicHqZH7Ku+ODWKjo6FI
QNTOM39uT6BAtMMrjESjuQxbpY52A5AefKsewwfBkROzLLMj2tK9U3whtrjY8nqW
fXkPnoUD9yFyROskT7Gt/EX6VJGq3AoG5VhefyDtg9W+khCHphF7KRgFAaiTdptl
NYtIabpOaAMY9U1r/qK1zX3A+q8BQBIB83RQ0OhHh1in1hJOtOox0wZwNjKVDmbO
h0n3N0VnGClNwOtlSaB4LYp7F+XYeNKJ/S/DtITrARHCv1pDaSZZInDhJFeODOqH
Eb75BDuSQiBe1Qcl+1KsnSMj9dvpgnkFuD8VzUU6Sd4FO8N5dLfybb2JKX0MOOT3
I5laxM1LmcpYxKmoUylxKhPjBlSsrNNlBRX90yIayKEEsYZHNnpv985IKP8Gf8Yj
KbVMUTW7oUl8XjbpjLCGmfvb0pmVI3r53UD8YriW7lFZdWj14xGr0daWJr7yuM6f
ewkGT8aNmofwGBbYA6qO7o7U2Fje8nq4bsLys2UhilqAwU49kAY765rs+UIHcp5+
PD/ZOPudEpsnBatqISNCsNFDR8gScS85HE4gFN4ddbEkto9gQFvkbEyfKlhz9fsQ
4WQm1RuOWw4CpxU4yQOnl8LrPNHe6IPFVkpoU6bv8+IODQWs3Qn99a2C8yCr89vS
BYdz6O1cWaPTCKujEnQI2/lpdi7Dy/KUjQLx3hltkEDyl7NKCM93o8n+FU8l2YDz
I6NXwVav8gw5owQMyAUJJ5EGD/6jRs46jaVWnIwZcWw48/OWBotCHnU5omtr6f2i
rwTGQ9qByHNbFcb13X2iv+ZOtnTqSPxVLz6TpAn3jamE6aeudIDX/V+Z0+ElOWru
UK4e9wYvGxAsdeE2RNhYUnH4wiOpRGXwLKxAY67p/TkAJs0ToSfgTO677reO2k21
UL0061ZZYbZX2OQdlUb9MaOMZkVUIpvoHpJfjCwOJ/dGF00G5mpL/3Tvg7wNgrxO
aElK7Pffocp7Yu6vCqfdXGkh0BZrb8ZmtERw18Ly5Bg2PSsI+8WblmaO6lk+Yk/F
Wt5rRd+jsnjrkx7s0EK9eGDhwGLOLT77iIREmqq1tx8vds5WDVcEulnwLqq9Pf2g
oHOQiyRAiaEYxhzBco6q30Cnf9IPkfnVeD6rad674GW7sO3HPwbg/R9wo4KF8+Zc
YDeLaSE3MgHzxkwehMa98DACOdeYpFwlEYSDyUujoTZ3cX0eKmfqcBPk3V96pd0d
d9rk7fWmKH7JUv0mVoitIFSjUd/9S9yBNU8n2mAQWT/vJtx1TOAbc5wqroVuT/P5
ZQvGv+cLPk1lX0t4LiNF3tlDx2ixrSnRmDHkDKedqKrQ4HZhXTv7+3WBVgrUGePV
BeAxXIe7ut9eOb48htvjuvDXiS9CibM3YzL6VPy1j9aYY5PtV+ihhBLfsv7tolea
CCLPtJpV6zO7K0t+zmM1fXiSm9mXu6hGeIBfSSvQ+ISft8FICPmymsKwfvJL3QMB
lLLG/sdWx3BtqLo1wP8MPI5J3Ig9ixQvECc2C+bwsKtu9+feY2wfJe5e2SXfjZDR
1mHdLbWFx3jdpRisPB9aDhQyVi1KN0Yb2f9mTRoXfD//aKaCqJG65Sd4AvQ8pJz7
x/TIfp+h2jaZ46yLXxzcPjUuAeav0xv5NQERg4qz/1Mptwt/KsE/8GEmIMDuIsKC
EMjaxzx/ldROmLl1Dki+NkLKdbKCh06Dgb7Z5mG3sslhSEghNYLnGhTVRaWagDeH
o5+TY7UOu3n0vU3M23PfNf+b+Ppb0IiwJGc2+xBVtgwMTf2Nn0Sv4Snu9GuJLLx3
wC/BfwECjp2i+ZLhVQEqwyhGB9Mcru6iZa5MghwVWJ+QcSQFiL6DeWAg8yJQi3LQ
RHJCMfcR9Ee2WOj5D+me9Rdh+M3DPml4dhXKV7cZs0h2Xe0sJy2JSXfinfmtL+9Z
YWt/Y3rowtIZ9qAT/8qXJY75U/nCSYQDj9N9mObdk9dNV3NfHuMEJ1PcvN+505EV
zG5qpZitOkaamMH5otBwy+GilDJhwur5MA7WoQOtjuv4zxqZVAHKD8dgJpdX9WZT
Tpu7VzK5Ax8KwQi6wZBAEzCDoU3yW04CEwEimqvU1iQECfDwK0w8A0wUYH4I2DAq
eUm4xzKHHlNTJoWgPRoPTEoeqKm8emxDbJ/0bhnUvlR7kIoRzOIVKUWTvY6v7gTW
Ey7NTD37K+U+4Rt+T6R+sOaIpIatXHMY7Olo9HJr/3XrxXKmf8umh86SdsZe6mR3
3S8AJDHORw8smdfHbbT8l+OLxISNBvEHKi3GXm1aVwhGw2CuDYs7b+xTwT7cl5tb
pjlondZj/i7F/zg6N9OSesFypCd9LvVGlhPAUTFtf+p3eG7sWXFeUx8NbI8SDh9j
MrfcjQyvL+Cc6liWbeyX1+JIULfJZu90niwoH4mq+XYN/6WjlKywM/JBVu24h5ii
WQFWLkuwqtI18Fh9LDeRSID/XLYbSL5SinaBJzLwCLyyChzipO2BQc9JnlIiRt80
mKS8SnkQ+ltIrOXLucJs3BoQBk3YxTM8QS4RSEvT0mhxGAh8rYIpkunh/VLEI2Xc
qyBKxZFwev31f2obSqzpJYr2+yhg5cDrSBmhemNcxfUN7HENNNstM8X/q7A1FWjO
8VqupzDdI3pWTAtJ2ZbyjrmrAdN9kYDLgmG++NI4mVNwv897TUcSTlrfMu9uCFkq
6Wnq/eNyXKeYZyfnRFBk0nT2x9P6dchEPRKxBgwMfxiy6EPBi/+BmTr5OpuKbNj4
0A4PHyHpwrFCrqudxklQBpR0ulhQ9GXHn4o2lxzzUPddf5d13T3dKW8S8X61rbNM
ClpW9kmjx/9cM1o+Nce+i2NDh4POq6ksz0t65zXjO5ZbU4+pDXV69WHQ/+YaJv26
qdRsTw2N8jEJGRurO55U7io9z6YcAtVFjyDi6bbLO4louDXFqKuqXhQHP7hITtxg
1+E1nYF1EI3j17m8+VQvZQXmPBXaMadEAvgERIzW+XgE5Q/1HZREZHvIv2r46j1F
mYR+oUEV44k+p7i1nJwtaM53zewiXlaz95YwjcaQvo/elSud/oNCyoP0Wr4+X7CZ
qGNh6TiI+ryxpvgIdFEhvFOlxIFpRQRRzWeBSZhiWLa18UJC0d4Gictu7LXnRiOF
USFTLF276qByAoH/zQSl452lJqJjedY3l2K6e/E4Z/AI/OmJsBWlDN02Uc8ubnah
oPre5iz5PLhU2+/Z3lJCDzqfhjkERqNvUCMU1pCKu6GmajDJtqiuU1dwkfo+0/0J
bU1DTCU5iOyJ2cTJ6lslXeyGKLq7uN5rOOj5Tb1LsAYTacBfKXOUab//acCaYRSV
bd8RsfR6EUcGeSnHpk1VD56v5QIhLelMkBcFlr0kAv1J67jbfqetbtsELuOhLEmp
sYPnftIdXVvuoF5OWj60ReBWFIlUe1Xm6UUr7iFbhwBewbZodJvr6/Cq9efSb8Lh
YCamKT1jrICYTjRdR3qyya+/ZHuUfcqEK9MCI7wzYG9M1hehjV4BxNJdXbOcuk7J
BoIHY54fa19Vm10Txg/9JZn6fiI47C/cTSrinNPsckra+QkPtTi8VUp4w14dM1Ps
`protect end_protected
